`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2024/01/06 18:16:08
// Design Name: 
// Module Name: outputpicture
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module outputpicture(
    input vga_clk,
    input [31:0]rabbitout,
    input [31:0]chickenout,
    input rst_n,
    input data_read_active,
    input picture_active,
    input [9:0]h_addr,
    input [9:0]v_addr,
    output reg[3:0]outputrdata,
    output reg[3:0]outputgdata,
    output reg[3:0]outputbdata
    );
    // reg [18:0]addr;
    // wire [3:0]data_romr1; data_romg1; data_romb1;
    // wire [3:0]data_romr2; data_romg2; data_romb2;
    // wire picture_exist1; picture_exist2;
    // wire data_require; data_require1; data_require2;
    // wire [24:0]rabbit_exist; rabbit_require;
    // wire [49:0]chicken_exist; chicken_require;
    parameter
    HEIGHT = 10'd55,
    WIDTH = 10'd55,
    RMAR = 10'd22,
    LMAR = 10'd23,
    MAR = 10'd5;


    reg [3:0]r_chickenpic[3024:0];
    reg [3:0]g_chickenpic[3024:0];
    reg [3:0]b_chickenpic[3024:0];
    reg [3:0]r_rabbitpic[3024:0];
    reg [3:0]g_rabbitpic[3024:0];
    reg [3:0]b_rabbitpic[3024:0];

    always @(posedge vga_clk) begin
        if(!rst_n) begin
            outputrdata <= 4'b0; outputgdata <= 4'b0; outputbdata <= 4'b0;
        end


        //***********************     row0     ***************************//
        
        else if (v_addr >= 0*(HEIGHT + MAR)  && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd0) begin   //(0;0)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd1) begin   //(0;1)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd2) begin   //(0;2)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd3) begin   //(0;3)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd4) begin   //(0;4)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd5) begin   //(0;5)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd6) begin   //(0;6)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd7) begin   //(0;7)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd8) begin   //(0;8)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr >= 0*(HEIGHT + MAR) && v_addr < HEIGHT + 0*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd9) begin   //(0;9)
            outputrdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 0*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row1     ***************************//

        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd10) begin   //(1;0)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd11) begin   //(1;1)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd12) begin   //(1;2)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd13) begin   //(1;3)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd14) begin   //(1;4)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd15) begin   //(1;5)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd16) begin   //(1;6)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd17) begin   //(1;7)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd18) begin   //(1;8)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 1*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 1*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd19) begin   //(1;9)
            outputrdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 1*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row2     ***************************//

        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd20) begin   //(2;0)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd21) begin   //(2;1)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd22) begin   //(2;2)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd23) begin   //(2;3)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd24) begin   //(2;4)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd25) begin   //(2;5)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd26) begin   //(2;6)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd27) begin   //(2;7)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd28) begin   //(2;8)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 2*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 2*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd29) begin   //(2;9)
            outputrdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 2*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end
        
        //***********************     row3     ***************************//

        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd30) begin   //(3;0)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd31) begin   //(3;1)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd32) begin   //(3;2)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd33) begin   //(3;3)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd34) begin   //(3;4)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd35) begin   //(3;5)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd36) begin   //(3;6)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd37) begin   //(3;7)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd38) begin   //(3;8)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 3*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 3*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd39) begin   //(3;9)
            outputrdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 3*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row4     ***************************//

        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd40) begin   //(4;0)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd41) begin   //(4;1)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd42) begin   //(4;2)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd43) begin   //(4;3)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd44) begin   //(4;4)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd45) begin   //(4;5)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd46) begin   //(4;6)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd47) begin   //(4;7)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd48) begin   //(4;8)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 4*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 4*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && rabbitout >= 32'd0 &&chickenout > 32'd49) begin   //(4;9)
            outputrdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_chickenpic[(v_addr - 4*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row5     ***************************//

        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd0) begin   //(5;0)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd1) begin   //(5;1)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd2) begin   //(5;2)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd3) begin   //(5;3)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd4) begin   //(5;4)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd5) begin   //(5;5)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd6) begin   //(5;6)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd7) begin   //(5;7)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd8) begin   //(5;8)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 5*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 5*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd9) begin   //(5;9)
            outputrdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 5*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row6     ***************************//

        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd10) begin   //(6;0)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd11) begin   //(6;1)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd12) begin   //(6;2)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd13) begin   //(6;3)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd14) begin   //(6;4)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 5*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 5*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd15) begin   //(6;5)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 5*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 6*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 6*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd16) begin   //(6;6)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 6*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 7*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 7*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd17) begin   //(6;7)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 7*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 8*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 8*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd18) begin   //(6;8)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 8*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 6*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 6*(HEIGHT + MAR) - 1 && h_addr > RMAR + 9*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 9*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd19) begin   //(6;9)
            outputrdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 6*(HEIGHT + MAR))*WIDTH + (h_addr - 9*(WIDTH + MAR) - RMAR)];
        end

        //***********************     row7     ***************************//

        else if (v_addr > 7*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 7*(HEIGHT + MAR) - 1 && h_addr > RMAR + 0*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 0*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd20) begin   //(7;0)
            outputrdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 0*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 7*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 7*(HEIGHT + MAR) - 1 && h_addr > RMAR + 1*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 1*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd21) begin   //(7;1)
            outputrdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 1*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 7*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 7*(HEIGHT + MAR) - 1 && h_addr > RMAR + 2*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 2*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd22) begin   //(7;2)
            outputrdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 2*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 7*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 7*(HEIGHT + MAR) - 1 && h_addr > RMAR + 3*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 3*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd23) begin   //(7;3)
            outputrdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 3*(WIDTH + MAR) - RMAR)];
        end
        else if (v_addr > 7*(HEIGHT + MAR) - 1 && v_addr < HEIGHT + 7*(HEIGHT + MAR) - 1 && h_addr > RMAR + 4*(WIDTH + MAR) - 1 && h_addr < RMAR + WIDTH + 4*(WIDTH + MAR) - 1 && chickenout < 32'd51 && rabbitout < 32'd26 && chickenout >= 32'd0  && rabbitout > 32'd24) begin   //(7;4)
            outputrdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputgdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
            outputbdata <= r_rabbitpic[(v_addr - 7*(HEIGHT + MAR))*WIDTH + (h_addr - 4*(WIDTH + MAR) - RMAR)];
        end
        else begin 
            outputrdata <= 4'b1111;
            outputgdata <= 4'b1111;
            outputbdata <= 4'b1111;
        end
    end

    always @(negedge rst_n) begin
        r_chickenpic[0] <= 4'b1111;
        r_chickenpic[1] <= 4'b1111;
        r_chickenpic[2] <= 4'b1111;
        r_chickenpic[3] <= 4'b1111;
        r_chickenpic[4] <= 4'b1111;
        r_chickenpic[5] <= 4'b1111;
        r_chickenpic[6] <= 4'b1111;
        r_chickenpic[7] <= 4'b1111;
        r_chickenpic[8] <= 4'b1111;
        r_chickenpic[9] <= 4'b1111;
        r_chickenpic[10] <= 4'b1111;
        r_chickenpic[11] <= 4'b1111;
        r_chickenpic[12] <= 4'b1111;
        r_chickenpic[13] <= 4'b1111;
        r_chickenpic[14] <= 4'b1111;
        r_chickenpic[15] <= 4'b1111;
        r_chickenpic[16] <= 4'b1111;
        r_chickenpic[17] <= 4'b1111;
        r_chickenpic[18] <= 4'b1111;
        r_chickenpic[19] <= 4'b1111;
        r_chickenpic[20] <= 4'b1111;
        r_chickenpic[21] <= 4'b1111;
        r_chickenpic[22] <= 4'b1111;
        r_chickenpic[23] <= 4'b1111;
        r_chickenpic[24] <= 4'b1111;
        r_chickenpic[25] <= 4'b1111;
        r_chickenpic[26] <= 4'b1111;
        r_chickenpic[27] <= 4'b1111;
        r_chickenpic[28] <= 4'b1111;
        r_chickenpic[29] <= 4'b1111;
        r_chickenpic[30] <= 4'b1111;
        r_chickenpic[31] <= 4'b1111;
        r_chickenpic[32] <= 4'b1111;
        r_chickenpic[33] <= 4'b1111;
        r_chickenpic[34] <= 4'b1111;
        r_chickenpic[35] <= 4'b1111;
        r_chickenpic[36] <= 4'b1111;
        r_chickenpic[37] <= 4'b1111;
        r_chickenpic[38] <= 4'b1111;
        r_chickenpic[39] <= 4'b1111;
        r_chickenpic[40] <= 4'b1111;
        r_chickenpic[41] <= 4'b1111;
        r_chickenpic[42] <= 4'b1111;
        r_chickenpic[43] <= 4'b1111;
        r_chickenpic[44] <= 4'b1111;
        r_chickenpic[45] <= 4'b1111;
        r_chickenpic[46] <= 4'b1111;
        r_chickenpic[47] <= 4'b1111;
        r_chickenpic[48] <= 4'b1111;
        r_chickenpic[49] <= 4'b1111;
        r_chickenpic[50] <= 4'b1111;
        r_chickenpic[51] <= 4'b1111;
        r_chickenpic[52] <= 4'b1111;
        r_chickenpic[53] <= 4'b1111;
        r_chickenpic[54] <= 4'b1111;
        r_chickenpic[55] <= 4'b1111;
        r_chickenpic[56] <= 4'b1111;
        r_chickenpic[57] <= 4'b1111;
        r_chickenpic[58] <= 4'b1111;
        r_chickenpic[59] <= 4'b1111;
        r_chickenpic[60] <= 4'b1111;
        r_chickenpic[61] <= 4'b1111;
        r_chickenpic[62] <= 4'b1111;
        r_chickenpic[63] <= 4'b1111;
        r_chickenpic[64] <= 4'b1111;
        r_chickenpic[65] <= 4'b1111;
        r_chickenpic[66] <= 4'b1111;
        r_chickenpic[67] <= 4'b1111;
        r_chickenpic[68] <= 4'b1111;
        r_chickenpic[69] <= 4'b1111;
        r_chickenpic[70] <= 4'b1111;
        r_chickenpic[71] <= 4'b1111;
        r_chickenpic[72] <= 4'b1111;
        r_chickenpic[73] <= 4'b1111;
        r_chickenpic[74] <= 4'b1111;
        r_chickenpic[75] <= 4'b1111;
        r_chickenpic[76] <= 4'b1111;
        r_chickenpic[77] <= 4'b1111;
        r_chickenpic[78] <= 4'b1111;
        r_chickenpic[79] <= 4'b1111;
        r_chickenpic[80] <= 4'b1111;
        r_chickenpic[81] <= 4'b1111;
        r_chickenpic[82] <= 4'b1111;
        r_chickenpic[83] <= 4'b1111;
        r_chickenpic[84] <= 4'b1111;
        r_chickenpic[85] <= 4'b1111;
        r_chickenpic[86] <= 4'b1111;
        r_chickenpic[87] <= 4'b1111;
        r_chickenpic[88] <= 4'b1111;
        r_chickenpic[89] <= 4'b1111;
        r_chickenpic[90] <= 4'b1111;
        r_chickenpic[91] <= 4'b1111;
        r_chickenpic[92] <= 4'b1111;
        r_chickenpic[93] <= 4'b1111;
        r_chickenpic[94] <= 4'b1111;
        r_chickenpic[95] <= 4'b1111;
        r_chickenpic[96] <= 4'b1111;
        r_chickenpic[97] <= 4'b1111;
        r_chickenpic[98] <= 4'b1111;
        r_chickenpic[99] <= 4'b1111;
        r_chickenpic[100] <= 4'b1111;
        r_chickenpic[101] <= 4'b1111;
        r_chickenpic[102] <= 4'b1111;
        r_chickenpic[103] <= 4'b1111;
        r_chickenpic[104] <= 4'b1111;
        r_chickenpic[105] <= 4'b1111;
        r_chickenpic[106] <= 4'b1111;
        r_chickenpic[107] <= 4'b1111;
        r_chickenpic[108] <= 4'b1111;
        r_chickenpic[109] <= 4'b1111;
        r_chickenpic[110] <= 4'b1111;
        r_chickenpic[111] <= 4'b1111;
        r_chickenpic[112] <= 4'b1111;
        r_chickenpic[113] <= 4'b1111;
        r_chickenpic[114] <= 4'b1111;
        r_chickenpic[115] <= 4'b1111;
        r_chickenpic[116] <= 4'b1111;
        r_chickenpic[117] <= 4'b1111;
        r_chickenpic[118] <= 4'b1111;
        r_chickenpic[119] <= 4'b1111;
        r_chickenpic[120] <= 4'b1111;
        r_chickenpic[121] <= 4'b1111;
        r_chickenpic[122] <= 4'b1111;
        r_chickenpic[123] <= 4'b1111;
        r_chickenpic[124] <= 4'b1111;
        r_chickenpic[125] <= 4'b1111;
        r_chickenpic[126] <= 4'b1111;
        r_chickenpic[127] <= 4'b1111;
        r_chickenpic[128] <= 4'b1111;
        r_chickenpic[129] <= 4'b1111;
        r_chickenpic[130] <= 4'b1111;
        r_chickenpic[131] <= 4'b1111;
        r_chickenpic[132] <= 4'b1111;
        r_chickenpic[133] <= 4'b1111;
        r_chickenpic[134] <= 4'b1111;
        r_chickenpic[135] <= 4'b1111;
        r_chickenpic[136] <= 4'b1111;
        r_chickenpic[137] <= 4'b1111;
        r_chickenpic[138] <= 4'b1111;
        r_chickenpic[139] <= 4'b1111;
        r_chickenpic[140] <= 4'b1111;
        r_chickenpic[141] <= 4'b1111;
        r_chickenpic[142] <= 4'b1111;
        r_chickenpic[143] <= 4'b1111;
        r_chickenpic[144] <= 4'b1111;
        r_chickenpic[145] <= 4'b1111;
        r_chickenpic[146] <= 4'b1111;
        r_chickenpic[147] <= 4'b1111;
        r_chickenpic[148] <= 4'b1111;
        r_chickenpic[149] <= 4'b1111;
        r_chickenpic[150] <= 4'b1111;
        r_chickenpic[151] <= 4'b1111;
        r_chickenpic[152] <= 4'b1111;
        r_chickenpic[153] <= 4'b1111;
        r_chickenpic[154] <= 4'b1111;
        r_chickenpic[155] <= 4'b1111;
        r_chickenpic[156] <= 4'b1111;
        r_chickenpic[157] <= 4'b1111;
        r_chickenpic[158] <= 4'b1111;
        r_chickenpic[159] <= 4'b1111;
        r_chickenpic[160] <= 4'b1111;
        r_chickenpic[161] <= 4'b1111;
        r_chickenpic[162] <= 4'b1111;
        r_chickenpic[163] <= 4'b1111;
        r_chickenpic[164] <= 4'b1111;
        r_chickenpic[165] <= 4'b1111;
        r_chickenpic[166] <= 4'b1111;
        r_chickenpic[167] <= 4'b1111;
        r_chickenpic[168] <= 4'b1111;
        r_chickenpic[169] <= 4'b1111;
        r_chickenpic[170] <= 4'b1111;
        r_chickenpic[171] <= 4'b1111;
        r_chickenpic[172] <= 4'b1111;
        r_chickenpic[173] <= 4'b1111;
        r_chickenpic[174] <= 4'b1111;
        r_chickenpic[175] <= 4'b1111;
        r_chickenpic[176] <= 4'b1111;
        r_chickenpic[177] <= 4'b1111;
        r_chickenpic[178] <= 4'b1111;
        r_chickenpic[179] <= 4'b1111;
        r_chickenpic[180] <= 4'b1111;
        r_chickenpic[181] <= 4'b1111;
        r_chickenpic[182] <= 4'b1111;
        r_chickenpic[183] <= 4'b1111;
        r_chickenpic[184] <= 4'b1111;
        r_chickenpic[185] <= 4'b1111;
        r_chickenpic[186] <= 4'b1111;
        r_chickenpic[187] <= 4'b1111;
        r_chickenpic[188] <= 4'b1111;
        r_chickenpic[189] <= 4'b1111;
        r_chickenpic[190] <= 4'b1111;
        r_chickenpic[191] <= 4'b1111;
        r_chickenpic[192] <= 4'b1111;
        r_chickenpic[193] <= 4'b1111;
        r_chickenpic[194] <= 4'b1111;
        r_chickenpic[195] <= 4'b1111;
        r_chickenpic[196] <= 4'b1111;
        r_chickenpic[197] <= 4'b1111;
        r_chickenpic[198] <= 4'b1111;
        r_chickenpic[199] <= 4'b1111;
        r_chickenpic[200] <= 4'b1111;
        r_chickenpic[201] <= 4'b1111;
        r_chickenpic[202] <= 4'b1111;
        r_chickenpic[203] <= 4'b1111;
        r_chickenpic[204] <= 4'b1111;
        r_chickenpic[205] <= 4'b1111;
        r_chickenpic[206] <= 4'b1111;
        r_chickenpic[207] <= 4'b1111;
        r_chickenpic[208] <= 4'b1111;
        r_chickenpic[209] <= 4'b1111;
        r_chickenpic[210] <= 4'b1111;
        r_chickenpic[211] <= 4'b1111;
        r_chickenpic[212] <= 4'b1111;
        r_chickenpic[213] <= 4'b1111;
        r_chickenpic[214] <= 4'b1111;
        r_chickenpic[215] <= 4'b1111;
        r_chickenpic[216] <= 4'b1111;
        r_chickenpic[217] <= 4'b1111;
        r_chickenpic[218] <= 4'b1111;
        r_chickenpic[219] <= 4'b1111;
        r_chickenpic[220] <= 4'b1111;
        r_chickenpic[221] <= 4'b1111;
        r_chickenpic[222] <= 4'b1111;
        r_chickenpic[223] <= 4'b1111;
        r_chickenpic[224] <= 4'b1111;
        r_chickenpic[225] <= 4'b1111;
        r_chickenpic[226] <= 4'b1111;
        r_chickenpic[227] <= 4'b1111;
        r_chickenpic[228] <= 4'b1111;
        r_chickenpic[229] <= 4'b1111;
        r_chickenpic[230] <= 4'b1111;
        r_chickenpic[231] <= 4'b1111;
        r_chickenpic[232] <= 4'b1111;
        r_chickenpic[233] <= 4'b1111;
        r_chickenpic[234] <= 4'b1111;
        r_chickenpic[235] <= 4'b1111;
        r_chickenpic[236] <= 4'b1111;
        r_chickenpic[237] <= 4'b1111;
        r_chickenpic[238] <= 4'b1111;
        r_chickenpic[239] <= 4'b1111;
        r_chickenpic[240] <= 4'b1111;
        r_chickenpic[241] <= 4'b1111;
        r_chickenpic[242] <= 4'b1111;
        r_chickenpic[243] <= 4'b1111;
        r_chickenpic[244] <= 4'b1111;
        r_chickenpic[245] <= 4'b1111;
        r_chickenpic[246] <= 4'b1111;
        r_chickenpic[247] <= 4'b1111;
        r_chickenpic[248] <= 4'b1111;
        r_chickenpic[249] <= 4'b1111;
        r_chickenpic[250] <= 4'b1111;
        r_chickenpic[251] <= 4'b1111;
        r_chickenpic[252] <= 4'b1111;
        r_chickenpic[253] <= 4'b1111;
        r_chickenpic[254] <= 4'b1111;
        r_chickenpic[255] <= 4'b1111;
        r_chickenpic[256] <= 4'b1111;
        r_chickenpic[257] <= 4'b1111;
        r_chickenpic[258] <= 4'b1111;
        r_chickenpic[259] <= 4'b1111;
        r_chickenpic[260] <= 4'b1111;
        r_chickenpic[261] <= 4'b1111;
        r_chickenpic[262] <= 4'b1111;
        r_chickenpic[263] <= 4'b1111;
        r_chickenpic[264] <= 4'b1111;
        r_chickenpic[265] <= 4'b1111;
        r_chickenpic[266] <= 4'b1111;
        r_chickenpic[267] <= 4'b1111;
        r_chickenpic[268] <= 4'b1111;
        r_chickenpic[269] <= 4'b1111;
        r_chickenpic[270] <= 4'b1111;
        r_chickenpic[271] <= 4'b1111;
        r_chickenpic[272] <= 4'b1111;
        r_chickenpic[273] <= 4'b1111;
        r_chickenpic[274] <= 4'b1111;
        r_chickenpic[275] <= 4'b1111;
        r_chickenpic[276] <= 4'b1111;
        r_chickenpic[277] <= 4'b1111;
        r_chickenpic[278] <= 4'b1111;
        r_chickenpic[279] <= 4'b1111;
        r_chickenpic[280] <= 4'b1111;
        r_chickenpic[281] <= 4'b1111;
        r_chickenpic[282] <= 4'b1111;
        r_chickenpic[283] <= 4'b1111;
        r_chickenpic[284] <= 4'b1111;
        r_chickenpic[285] <= 4'b1111;
        r_chickenpic[286] <= 4'b1111;
        r_chickenpic[287] <= 4'b1111;
        r_chickenpic[288] <= 4'b1111;
        r_chickenpic[289] <= 4'b1111;
        r_chickenpic[290] <= 4'b1111;
        r_chickenpic[291] <= 4'b1111;
        r_chickenpic[292] <= 4'b1111;
        r_chickenpic[293] <= 4'b1111;
        r_chickenpic[294] <= 4'b1111;
        r_chickenpic[295] <= 4'b1111;
        r_chickenpic[296] <= 4'b1111;
        r_chickenpic[297] <= 4'b1111;
        r_chickenpic[298] <= 4'b1111;
        r_chickenpic[299] <= 4'b1111;
        r_chickenpic[300] <= 4'b0000;
        r_chickenpic[301] <= 4'b0000;
        r_chickenpic[302] <= 4'b1111;
        r_chickenpic[303] <= 4'b1111;
        r_chickenpic[304] <= 4'b1111;
        r_chickenpic[305] <= 4'b1111;
        r_chickenpic[306] <= 4'b1111;
        r_chickenpic[307] <= 4'b1111;
        r_chickenpic[308] <= 4'b1111;
        r_chickenpic[309] <= 4'b1111;
        r_chickenpic[310] <= 4'b1111;
        r_chickenpic[311] <= 4'b1111;
        r_chickenpic[312] <= 4'b1111;
        r_chickenpic[313] <= 4'b1111;
        r_chickenpic[314] <= 4'b1111;
        r_chickenpic[315] <= 4'b1111;
        r_chickenpic[316] <= 4'b1111;
        r_chickenpic[317] <= 4'b1111;
        r_chickenpic[318] <= 4'b1111;
        r_chickenpic[319] <= 4'b1111;
        r_chickenpic[320] <= 4'b1111;
        r_chickenpic[321] <= 4'b1111;
        r_chickenpic[322] <= 4'b1111;
        r_chickenpic[323] <= 4'b1111;
        r_chickenpic[324] <= 4'b1111;
        r_chickenpic[325] <= 4'b1111;
        r_chickenpic[326] <= 4'b1111;
        r_chickenpic[327] <= 4'b1111;
        r_chickenpic[328] <= 4'b1111;
        r_chickenpic[329] <= 4'b1111;
        r_chickenpic[330] <= 4'b1111;
        r_chickenpic[331] <= 4'b1111;
        r_chickenpic[332] <= 4'b1111;
        r_chickenpic[333] <= 4'b1111;
        r_chickenpic[334] <= 4'b1111;
        r_chickenpic[335] <= 4'b1111;
        r_chickenpic[336] <= 4'b1111;
        r_chickenpic[337] <= 4'b1111;
        r_chickenpic[338] <= 4'b1111;
        r_chickenpic[339] <= 4'b1111;
        r_chickenpic[340] <= 4'b1111;
        r_chickenpic[341] <= 4'b1111;
        r_chickenpic[342] <= 4'b1111;
        r_chickenpic[343] <= 4'b1111;
        r_chickenpic[344] <= 4'b1111;
        r_chickenpic[345] <= 4'b1111;
        r_chickenpic[346] <= 4'b1111;
        r_chickenpic[347] <= 4'b1111;
        r_chickenpic[348] <= 4'b1111;
        r_chickenpic[349] <= 4'b1111;
        r_chickenpic[350] <= 4'b1111;
        r_chickenpic[351] <= 4'b1111;
        r_chickenpic[352] <= 4'b1111;
        r_chickenpic[353] <= 4'b1111;
        r_chickenpic[354] <= 4'b0000;
        r_chickenpic[355] <= 4'b0000;
        r_chickenpic[356] <= 4'b0000;
        r_chickenpic[357] <= 4'b1111;
        r_chickenpic[358] <= 4'b1111;
        r_chickenpic[359] <= 4'b1111;
        r_chickenpic[360] <= 4'b1111;
        r_chickenpic[361] <= 4'b1111;
        r_chickenpic[362] <= 4'b1111;
        r_chickenpic[363] <= 4'b1111;
        r_chickenpic[364] <= 4'b1111;
        r_chickenpic[365] <= 4'b1111;
        r_chickenpic[366] <= 4'b1111;
        r_chickenpic[367] <= 4'b1111;
        r_chickenpic[368] <= 4'b1111;
        r_chickenpic[369] <= 4'b1111;
        r_chickenpic[370] <= 4'b1111;
        r_chickenpic[371] <= 4'b1111;
        r_chickenpic[372] <= 4'b1111;
        r_chickenpic[373] <= 4'b1111;
        r_chickenpic[374] <= 4'b1111;
        r_chickenpic[375] <= 4'b1111;
        r_chickenpic[376] <= 4'b1111;
        r_chickenpic[377] <= 4'b1111;
        r_chickenpic[378] <= 4'b1111;
        r_chickenpic[379] <= 4'b1111;
        r_chickenpic[380] <= 4'b1111;
        r_chickenpic[381] <= 4'b1111;
        r_chickenpic[382] <= 4'b1111;
        r_chickenpic[383] <= 4'b1111;
        r_chickenpic[384] <= 4'b1111;
        r_chickenpic[385] <= 4'b1111;
        r_chickenpic[386] <= 4'b1111;
        r_chickenpic[387] <= 4'b1111;
        r_chickenpic[388] <= 4'b1111;
        r_chickenpic[389] <= 4'b1111;
        r_chickenpic[390] <= 4'b1111;
        r_chickenpic[391] <= 4'b1111;
        r_chickenpic[392] <= 4'b1111;
        r_chickenpic[393] <= 4'b1111;
        r_chickenpic[394] <= 4'b1111;
        r_chickenpic[395] <= 4'b1111;
        r_chickenpic[396] <= 4'b1111;
        r_chickenpic[397] <= 4'b1111;
        r_chickenpic[398] <= 4'b1111;
        r_chickenpic[399] <= 4'b1111;
        r_chickenpic[400] <= 4'b1111;
        r_chickenpic[401] <= 4'b1111;
        r_chickenpic[402] <= 4'b1111;
        r_chickenpic[403] <= 4'b1111;
        r_chickenpic[404] <= 4'b1111;
        r_chickenpic[405] <= 4'b1111;
        r_chickenpic[406] <= 4'b1111;
        r_chickenpic[407] <= 4'b1111;
        r_chickenpic[408] <= 4'b0000;
        r_chickenpic[409] <= 4'b0000;
        r_chickenpic[410] <= 4'b0000;
        r_chickenpic[411] <= 4'b0000;
        r_chickenpic[412] <= 4'b1111;
        r_chickenpic[413] <= 4'b1111;
        r_chickenpic[414] <= 4'b1111;
        r_chickenpic[415] <= 4'b1111;
        r_chickenpic[416] <= 4'b1111;
        r_chickenpic[417] <= 4'b1111;
        r_chickenpic[418] <= 4'b1111;
        r_chickenpic[419] <= 4'b1111;
        r_chickenpic[420] <= 4'b1111;
        r_chickenpic[421] <= 4'b1111;
        r_chickenpic[422] <= 4'b1111;
        r_chickenpic[423] <= 4'b1111;
        r_chickenpic[424] <= 4'b1111;
        r_chickenpic[425] <= 4'b1111;
        r_chickenpic[426] <= 4'b1111;
        r_chickenpic[427] <= 4'b1111;
        r_chickenpic[428] <= 4'b1111;
        r_chickenpic[429] <= 4'b1111;
        r_chickenpic[430] <= 4'b1111;
        r_chickenpic[431] <= 4'b1111;
        r_chickenpic[432] <= 4'b1111;
        r_chickenpic[433] <= 4'b1111;
        r_chickenpic[434] <= 4'b1111;
        r_chickenpic[435] <= 4'b1111;
        r_chickenpic[436] <= 4'b1111;
        r_chickenpic[437] <= 4'b1111;
        r_chickenpic[438] <= 4'b1111;
        r_chickenpic[439] <= 4'b1111;
        r_chickenpic[440] <= 4'b1111;
        r_chickenpic[441] <= 4'b1111;
        r_chickenpic[442] <= 4'b1111;
        r_chickenpic[443] <= 4'b1111;
        r_chickenpic[444] <= 4'b1111;
        r_chickenpic[445] <= 4'b1111;
        r_chickenpic[446] <= 4'b1111;
        r_chickenpic[447] <= 4'b1111;
        r_chickenpic[448] <= 4'b1111;
        r_chickenpic[449] <= 4'b1111;
        r_chickenpic[450] <= 4'b1111;
        r_chickenpic[451] <= 4'b1111;
        r_chickenpic[452] <= 4'b1111;
        r_chickenpic[453] <= 4'b1111;
        r_chickenpic[454] <= 4'b1111;
        r_chickenpic[455] <= 4'b1111;
        r_chickenpic[456] <= 4'b1111;
        r_chickenpic[457] <= 4'b1111;
        r_chickenpic[458] <= 4'b1111;
        r_chickenpic[459] <= 4'b1111;
        r_chickenpic[460] <= 4'b1111;
        r_chickenpic[461] <= 4'b1111;
        r_chickenpic[462] <= 4'b0000;
        r_chickenpic[463] <= 4'b0000;
        r_chickenpic[464] <= 4'b1111;
        r_chickenpic[465] <= 4'b0000;
        r_chickenpic[466] <= 4'b0000;
        r_chickenpic[467] <= 4'b1111;
        r_chickenpic[468] <= 4'b1111;
        r_chickenpic[469] <= 4'b1111;
        r_chickenpic[470] <= 4'b1111;
        r_chickenpic[471] <= 4'b1111;
        r_chickenpic[472] <= 4'b1111;
        r_chickenpic[473] <= 4'b1111;
        r_chickenpic[474] <= 4'b1111;
        r_chickenpic[475] <= 4'b1111;
        r_chickenpic[476] <= 4'b1111;
        r_chickenpic[477] <= 4'b1111;
        r_chickenpic[478] <= 4'b1111;
        r_chickenpic[479] <= 4'b1111;
        r_chickenpic[480] <= 4'b1111;
        r_chickenpic[481] <= 4'b1111;
        r_chickenpic[482] <= 4'b1111;
        r_chickenpic[483] <= 4'b1111;
        r_chickenpic[484] <= 4'b1111;
        r_chickenpic[485] <= 4'b1111;
        r_chickenpic[486] <= 4'b1111;
        r_chickenpic[487] <= 4'b1111;
        r_chickenpic[488] <= 4'b1111;
        r_chickenpic[489] <= 4'b1111;
        r_chickenpic[490] <= 4'b1111;
        r_chickenpic[491] <= 4'b1111;
        r_chickenpic[492] <= 4'b1111;
        r_chickenpic[493] <= 4'b1111;
        r_chickenpic[494] <= 4'b1111;
        r_chickenpic[495] <= 4'b1111;
        r_chickenpic[496] <= 4'b1111;
        r_chickenpic[497] <= 4'b1111;
        r_chickenpic[498] <= 4'b1111;
        r_chickenpic[499] <= 4'b1111;
        r_chickenpic[500] <= 4'b1111;
        r_chickenpic[501] <= 4'b1111;
        r_chickenpic[502] <= 4'b1111;
        r_chickenpic[503] <= 4'b1111;
        r_chickenpic[504] <= 4'b1111;
        r_chickenpic[505] <= 4'b1111;
        r_chickenpic[506] <= 4'b1111;
        r_chickenpic[507] <= 4'b1111;
        r_chickenpic[508] <= 4'b1111;
        r_chickenpic[509] <= 4'b1111;
        r_chickenpic[510] <= 4'b1111;
        r_chickenpic[511] <= 4'b1111;
        r_chickenpic[512] <= 4'b1111;
        r_chickenpic[513] <= 4'b0000;
        r_chickenpic[514] <= 4'b0000;
        r_chickenpic[515] <= 4'b0000;
        r_chickenpic[516] <= 4'b0000;
        r_chickenpic[517] <= 4'b0000;
        r_chickenpic[518] <= 4'b0000;
        r_chickenpic[519] <= 4'b1111;
        r_chickenpic[520] <= 4'b0000;
        r_chickenpic[521] <= 4'b0000;
        r_chickenpic[522] <= 4'b0000;
        r_chickenpic[523] <= 4'b0000;
        r_chickenpic[524] <= 4'b0000;
        r_chickenpic[525] <= 4'b0000;
        r_chickenpic[526] <= 4'b1111;
        r_chickenpic[527] <= 4'b1111;
        r_chickenpic[528] <= 4'b1111;
        r_chickenpic[529] <= 4'b1111;
        r_chickenpic[530] <= 4'b1111;
        r_chickenpic[531] <= 4'b1111;
        r_chickenpic[532] <= 4'b1111;
        r_chickenpic[533] <= 4'b1111;
        r_chickenpic[534] <= 4'b1111;
        r_chickenpic[535] <= 4'b1111;
        r_chickenpic[536] <= 4'b1111;
        r_chickenpic[537] <= 4'b1111;
        r_chickenpic[538] <= 4'b1111;
        r_chickenpic[539] <= 4'b1111;
        r_chickenpic[540] <= 4'b1111;
        r_chickenpic[541] <= 4'b1111;
        r_chickenpic[542] <= 4'b1111;
        r_chickenpic[543] <= 4'b1111;
        r_chickenpic[544] <= 4'b1111;
        r_chickenpic[545] <= 4'b1111;
        r_chickenpic[546] <= 4'b1111;
        r_chickenpic[547] <= 4'b1111;
        r_chickenpic[548] <= 4'b1111;
        r_chickenpic[549] <= 4'b1111;
        r_chickenpic[550] <= 4'b1111;
        r_chickenpic[551] <= 4'b1111;
        r_chickenpic[552] <= 4'b1111;
        r_chickenpic[553] <= 4'b1111;
        r_chickenpic[554] <= 4'b1111;
        r_chickenpic[555] <= 4'b1111;
        r_chickenpic[556] <= 4'b1111;
        r_chickenpic[557] <= 4'b1111;
        r_chickenpic[558] <= 4'b1111;
        r_chickenpic[559] <= 4'b1111;
        r_chickenpic[560] <= 4'b1111;
        r_chickenpic[561] <= 4'b1111;
        r_chickenpic[562] <= 4'b1111;
        r_chickenpic[563] <= 4'b1111;
        r_chickenpic[564] <= 4'b1111;
        r_chickenpic[565] <= 4'b0000;
        r_chickenpic[566] <= 4'b0000;
        r_chickenpic[567] <= 4'b0000;
        r_chickenpic[568] <= 4'b0000;
        r_chickenpic[569] <= 4'b0000;
        r_chickenpic[570] <= 4'b0000;
        r_chickenpic[571] <= 4'b0000;
        r_chickenpic[572] <= 4'b0000;
        r_chickenpic[573] <= 4'b0000;
        r_chickenpic[574] <= 4'b0000;
        r_chickenpic[575] <= 4'b0000;
        r_chickenpic[576] <= 4'b0000;
        r_chickenpic[577] <= 4'b0000;
        r_chickenpic[578] <= 4'b0000;
        r_chickenpic[579] <= 4'b0000;
        r_chickenpic[580] <= 4'b1111;
        r_chickenpic[581] <= 4'b1111;
        r_chickenpic[582] <= 4'b1111;
        r_chickenpic[583] <= 4'b1111;
        r_chickenpic[584] <= 4'b1111;
        r_chickenpic[585] <= 4'b1111;
        r_chickenpic[586] <= 4'b1111;
        r_chickenpic[587] <= 4'b1111;
        r_chickenpic[588] <= 4'b1111;
        r_chickenpic[589] <= 4'b1111;
        r_chickenpic[590] <= 4'b1111;
        r_chickenpic[591] <= 4'b1111;
        r_chickenpic[592] <= 4'b1111;
        r_chickenpic[593] <= 4'b1111;
        r_chickenpic[594] <= 4'b1111;
        r_chickenpic[595] <= 4'b1111;
        r_chickenpic[596] <= 4'b1111;
        r_chickenpic[597] <= 4'b1111;
        r_chickenpic[598] <= 4'b1111;
        r_chickenpic[599] <= 4'b1111;
        r_chickenpic[600] <= 4'b1111;
        r_chickenpic[601] <= 4'b1111;
        r_chickenpic[602] <= 4'b1111;
        r_chickenpic[603] <= 4'b1111;
        r_chickenpic[604] <= 4'b1111;
        r_chickenpic[605] <= 4'b1111;
        r_chickenpic[606] <= 4'b1111;
        r_chickenpic[607] <= 4'b1111;
        r_chickenpic[608] <= 4'b1111;
        r_chickenpic[609] <= 4'b1111;
        r_chickenpic[610] <= 4'b1111;
        r_chickenpic[611] <= 4'b1111;
        r_chickenpic[612] <= 4'b1111;
        r_chickenpic[613] <= 4'b1111;
        r_chickenpic[614] <= 4'b1111;
        r_chickenpic[615] <= 4'b1111;
        r_chickenpic[616] <= 4'b1111;
        r_chickenpic[617] <= 4'b1111;
        r_chickenpic[618] <= 4'b0000;
        r_chickenpic[619] <= 4'b0000;
        r_chickenpic[620] <= 4'b0000;
        r_chickenpic[621] <= 4'b1111;
        r_chickenpic[622] <= 4'b1111;
        r_chickenpic[623] <= 4'b1111;
        r_chickenpic[624] <= 4'b1111;
        r_chickenpic[625] <= 4'b1111;
        r_chickenpic[626] <= 4'b1111;
        r_chickenpic[627] <= 4'b1111;
        r_chickenpic[628] <= 4'b0000;
        r_chickenpic[629] <= 4'b0000;
        r_chickenpic[630] <= 4'b0000;
        r_chickenpic[631] <= 4'b1111;
        r_chickenpic[632] <= 4'b0000;
        r_chickenpic[633] <= 4'b0000;
        r_chickenpic[634] <= 4'b1111;
        r_chickenpic[635] <= 4'b1111;
        r_chickenpic[636] <= 4'b1111;
        r_chickenpic[637] <= 4'b1111;
        r_chickenpic[638] <= 4'b1111;
        r_chickenpic[639] <= 4'b1111;
        r_chickenpic[640] <= 4'b1111;
        r_chickenpic[641] <= 4'b1111;
        r_chickenpic[642] <= 4'b1111;
        r_chickenpic[643] <= 4'b1111;
        r_chickenpic[644] <= 4'b1111;
        r_chickenpic[645] <= 4'b1111;
        r_chickenpic[646] <= 4'b1111;
        r_chickenpic[647] <= 4'b1111;
        r_chickenpic[648] <= 4'b1111;
        r_chickenpic[649] <= 4'b1111;
        r_chickenpic[650] <= 4'b1111;
        r_chickenpic[651] <= 4'b1111;
        r_chickenpic[652] <= 4'b1111;
        r_chickenpic[653] <= 4'b1111;
        r_chickenpic[654] <= 4'b1111;
        r_chickenpic[655] <= 4'b1111;
        r_chickenpic[656] <= 4'b1111;
        r_chickenpic[657] <= 4'b1111;
        r_chickenpic[658] <= 4'b1111;
        r_chickenpic[659] <= 4'b1111;
        r_chickenpic[660] <= 4'b1111;
        r_chickenpic[661] <= 4'b1111;
        r_chickenpic[662] <= 4'b1111;
        r_chickenpic[663] <= 4'b1111;
        r_chickenpic[664] <= 4'b1111;
        r_chickenpic[665] <= 4'b1111;
        r_chickenpic[666] <= 4'b1111;
        r_chickenpic[667] <= 4'b1111;
        r_chickenpic[668] <= 4'b1111;
        r_chickenpic[669] <= 4'b1111;
        r_chickenpic[670] <= 4'b1111;
        r_chickenpic[671] <= 4'b1111;
        r_chickenpic[672] <= 4'b0000;
        r_chickenpic[673] <= 4'b0000;
        r_chickenpic[674] <= 4'b1111;
        r_chickenpic[675] <= 4'b1111;
        r_chickenpic[676] <= 4'b1111;
        r_chickenpic[677] <= 4'b1111;
        r_chickenpic[678] <= 4'b1111;
        r_chickenpic[679] <= 4'b1111;
        r_chickenpic[680] <= 4'b1111;
        r_chickenpic[681] <= 4'b1111;
        r_chickenpic[682] <= 4'b1111;
        r_chickenpic[683] <= 4'b1111;
        r_chickenpic[684] <= 4'b1111;
        r_chickenpic[685] <= 4'b0000;
        r_chickenpic[686] <= 4'b0000;
        r_chickenpic[687] <= 4'b0000;
        r_chickenpic[688] <= 4'b1111;
        r_chickenpic[689] <= 4'b1111;
        r_chickenpic[690] <= 4'b1111;
        r_chickenpic[691] <= 4'b1111;
        r_chickenpic[692] <= 4'b1111;
        r_chickenpic[693] <= 4'b1111;
        r_chickenpic[694] <= 4'b1111;
        r_chickenpic[695] <= 4'b1111;
        r_chickenpic[696] <= 4'b1111;
        r_chickenpic[697] <= 4'b1111;
        r_chickenpic[698] <= 4'b1111;
        r_chickenpic[699] <= 4'b1111;
        r_chickenpic[700] <= 4'b1111;
        r_chickenpic[701] <= 4'b1111;
        r_chickenpic[702] <= 4'b1111;
        r_chickenpic[703] <= 4'b1111;
        r_chickenpic[704] <= 4'b1111;
        r_chickenpic[705] <= 4'b1111;
        r_chickenpic[706] <= 4'b1111;
        r_chickenpic[707] <= 4'b1111;
        r_chickenpic[708] <= 4'b1111;
        r_chickenpic[709] <= 4'b1111;
        r_chickenpic[710] <= 4'b1111;
        r_chickenpic[711] <= 4'b1111;
        r_chickenpic[712] <= 4'b1111;
        r_chickenpic[713] <= 4'b1111;
        r_chickenpic[714] <= 4'b1111;
        r_chickenpic[715] <= 4'b1111;
        r_chickenpic[716] <= 4'b1111;
        r_chickenpic[717] <= 4'b1111;
        r_chickenpic[718] <= 4'b1111;
        r_chickenpic[719] <= 4'b1111;
        r_chickenpic[720] <= 4'b1111;
        r_chickenpic[721] <= 4'b1111;
        r_chickenpic[722] <= 4'b1111;
        r_chickenpic[723] <= 4'b1111;
        r_chickenpic[724] <= 4'b1111;
        r_chickenpic[725] <= 4'b1111;
        r_chickenpic[726] <= 4'b0000;
        r_chickenpic[727] <= 4'b0000;
        r_chickenpic[728] <= 4'b1111;
        r_chickenpic[729] <= 4'b1111;
        r_chickenpic[730] <= 4'b1111;
        r_chickenpic[731] <= 4'b1111;
        r_chickenpic[732] <= 4'b1111;
        r_chickenpic[733] <= 4'b0000;
        r_chickenpic[734] <= 4'b0000;
        r_chickenpic[735] <= 4'b0000;
        r_chickenpic[736] <= 4'b0000;
        r_chickenpic[737] <= 4'b1111;
        r_chickenpic[738] <= 4'b1111;
        r_chickenpic[739] <= 4'b1111;
        r_chickenpic[740] <= 4'b1111;
        r_chickenpic[741] <= 4'b0000;
        r_chickenpic[742] <= 4'b0000;
        r_chickenpic[743] <= 4'b1111;
        r_chickenpic[744] <= 4'b1111;
        r_chickenpic[745] <= 4'b1111;
        r_chickenpic[746] <= 4'b1111;
        r_chickenpic[747] <= 4'b1111;
        r_chickenpic[748] <= 4'b1111;
        r_chickenpic[749] <= 4'b1111;
        r_chickenpic[750] <= 4'b1111;
        r_chickenpic[751] <= 4'b1111;
        r_chickenpic[752] <= 4'b1111;
        r_chickenpic[753] <= 4'b1111;
        r_chickenpic[754] <= 4'b1111;
        r_chickenpic[755] <= 4'b1111;
        r_chickenpic[756] <= 4'b1111;
        r_chickenpic[757] <= 4'b1111;
        r_chickenpic[758] <= 4'b1111;
        r_chickenpic[759] <= 4'b1111;
        r_chickenpic[760] <= 4'b1111;
        r_chickenpic[761] <= 4'b1111;
        r_chickenpic[762] <= 4'b1111;
        r_chickenpic[763] <= 4'b1111;
        r_chickenpic[764] <= 4'b1111;
        r_chickenpic[765] <= 4'b1111;
        r_chickenpic[766] <= 4'b1111;
        r_chickenpic[767] <= 4'b1111;
        r_chickenpic[768] <= 4'b1111;
        r_chickenpic[769] <= 4'b1111;
        r_chickenpic[770] <= 4'b1111;
        r_chickenpic[771] <= 4'b1111;
        r_chickenpic[772] <= 4'b1111;
        r_chickenpic[773] <= 4'b1111;
        r_chickenpic[774] <= 4'b1111;
        r_chickenpic[775] <= 4'b1111;
        r_chickenpic[776] <= 4'b1111;
        r_chickenpic[777] <= 4'b1111;
        r_chickenpic[778] <= 4'b1111;
        r_chickenpic[779] <= 4'b1111;
        r_chickenpic[780] <= 4'b0000;
        r_chickenpic[781] <= 4'b0000;
        r_chickenpic[782] <= 4'b1111;
        r_chickenpic[783] <= 4'b1111;
        r_chickenpic[784] <= 4'b1111;
        r_chickenpic[785] <= 4'b1111;
        r_chickenpic[786] <= 4'b1111;
        r_chickenpic[787] <= 4'b1111;
        r_chickenpic[788] <= 4'b0000;
        r_chickenpic[789] <= 4'b0000;
        r_chickenpic[790] <= 4'b0000;
        r_chickenpic[791] <= 4'b0000;
        r_chickenpic[792] <= 4'b1111;
        r_chickenpic[793] <= 4'b1111;
        r_chickenpic[794] <= 4'b1111;
        r_chickenpic[795] <= 4'b1111;
        r_chickenpic[796] <= 4'b1111;
        r_chickenpic[797] <= 4'b0000;
        r_chickenpic[798] <= 4'b1111;
        r_chickenpic[799] <= 4'b1111;
        r_chickenpic[800] <= 4'b1111;
        r_chickenpic[801] <= 4'b1111;
        r_chickenpic[802] <= 4'b1111;
        r_chickenpic[803] <= 4'b1111;
        r_chickenpic[804] <= 4'b1111;
        r_chickenpic[805] <= 4'b1111;
        r_chickenpic[806] <= 4'b1111;
        r_chickenpic[807] <= 4'b1111;
        r_chickenpic[808] <= 4'b1111;
        r_chickenpic[809] <= 4'b1111;
        r_chickenpic[810] <= 4'b1111;
        r_chickenpic[811] <= 4'b1111;
        r_chickenpic[812] <= 4'b0000;
        r_chickenpic[813] <= 4'b0000;
        r_chickenpic[814] <= 4'b0000;
        r_chickenpic[815] <= 4'b1111;
        r_chickenpic[816] <= 4'b1111;
        r_chickenpic[817] <= 4'b1111;
        r_chickenpic[818] <= 4'b1111;
        r_chickenpic[819] <= 4'b1111;
        r_chickenpic[820] <= 4'b1111;
        r_chickenpic[821] <= 4'b1111;
        r_chickenpic[822] <= 4'b1111;
        r_chickenpic[823] <= 4'b1111;
        r_chickenpic[824] <= 4'b1111;
        r_chickenpic[825] <= 4'b1111;
        r_chickenpic[826] <= 4'b1111;
        r_chickenpic[827] <= 4'b1111;
        r_chickenpic[828] <= 4'b1111;
        r_chickenpic[829] <= 4'b1111;
        r_chickenpic[830] <= 4'b1111;
        r_chickenpic[831] <= 4'b1111;
        r_chickenpic[832] <= 4'b1111;
        r_chickenpic[833] <= 4'b1111;
        r_chickenpic[834] <= 4'b1111;
        r_chickenpic[835] <= 4'b0000;
        r_chickenpic[836] <= 4'b0000;
        r_chickenpic[837] <= 4'b1111;
        r_chickenpic[838] <= 4'b1111;
        r_chickenpic[839] <= 4'b1111;
        r_chickenpic[840] <= 4'b1111;
        r_chickenpic[841] <= 4'b1111;
        r_chickenpic[842] <= 4'b1111;
        r_chickenpic[843] <= 4'b0000;
        r_chickenpic[844] <= 4'b0000;
        r_chickenpic[845] <= 4'b0000;
        r_chickenpic[846] <= 4'b0000;
        r_chickenpic[847] <= 4'b1111;
        r_chickenpic[848] <= 4'b1111;
        r_chickenpic[849] <= 4'b1111;
        r_chickenpic[850] <= 4'b1111;
        r_chickenpic[851] <= 4'b1111;
        r_chickenpic[852] <= 4'b0000;
        r_chickenpic[853] <= 4'b0000;
        r_chickenpic[854] <= 4'b1111;
        r_chickenpic[855] <= 4'b1111;
        r_chickenpic[856] <= 4'b1111;
        r_chickenpic[857] <= 4'b1111;
        r_chickenpic[858] <= 4'b1111;
        r_chickenpic[859] <= 4'b1111;
        r_chickenpic[860] <= 4'b1111;
        r_chickenpic[861] <= 4'b1111;
        r_chickenpic[862] <= 4'b1111;
        r_chickenpic[863] <= 4'b1111;
        r_chickenpic[864] <= 4'b1111;
        r_chickenpic[865] <= 4'b0000;
        r_chickenpic[866] <= 4'b0000;
        r_chickenpic[867] <= 4'b0000;
        r_chickenpic[868] <= 4'b0000;
        r_chickenpic[869] <= 4'b0000;
        r_chickenpic[870] <= 4'b0000;
        r_chickenpic[871] <= 4'b1111;
        r_chickenpic[872] <= 4'b1111;
        r_chickenpic[873] <= 4'b1111;
        r_chickenpic[874] <= 4'b1111;
        r_chickenpic[875] <= 4'b1111;
        r_chickenpic[876] <= 4'b1111;
        r_chickenpic[877] <= 4'b1111;
        r_chickenpic[878] <= 4'b1111;
        r_chickenpic[879] <= 4'b1111;
        r_chickenpic[880] <= 4'b1111;
        r_chickenpic[881] <= 4'b1111;
        r_chickenpic[882] <= 4'b1111;
        r_chickenpic[883] <= 4'b1111;
        r_chickenpic[884] <= 4'b1111;
        r_chickenpic[885] <= 4'b1111;
        r_chickenpic[886] <= 4'b1111;
        r_chickenpic[887] <= 4'b1111;
        r_chickenpic[888] <= 4'b1111;
        r_chickenpic[889] <= 4'b0000;
        r_chickenpic[890] <= 4'b0000;
        r_chickenpic[891] <= 4'b1111;
        r_chickenpic[892] <= 4'b1111;
        r_chickenpic[893] <= 4'b1111;
        r_chickenpic[894] <= 4'b1111;
        r_chickenpic[895] <= 4'b1111;
        r_chickenpic[896] <= 4'b1111;
        r_chickenpic[897] <= 4'b1111;
        r_chickenpic[898] <= 4'b0000;
        r_chickenpic[899] <= 4'b0000;
        r_chickenpic[900] <= 4'b0000;
        r_chickenpic[901] <= 4'b0000;
        r_chickenpic[902] <= 4'b1111;
        r_chickenpic[903] <= 4'b1111;
        r_chickenpic[904] <= 4'b1111;
        r_chickenpic[905] <= 4'b1111;
        r_chickenpic[906] <= 4'b1111;
        r_chickenpic[907] <= 4'b0000;
        r_chickenpic[908] <= 4'b0000;
        r_chickenpic[909] <= 4'b1111;
        r_chickenpic[910] <= 4'b1111;
        r_chickenpic[911] <= 4'b1111;
        r_chickenpic[912] <= 4'b1111;
        r_chickenpic[913] <= 4'b1111;
        r_chickenpic[914] <= 4'b1111;
        r_chickenpic[915] <= 4'b1111;
        r_chickenpic[916] <= 4'b1111;
        r_chickenpic[917] <= 4'b1111;
        r_chickenpic[918] <= 4'b1111;
        r_chickenpic[919] <= 4'b0000;
        r_chickenpic[920] <= 4'b0000;
        r_chickenpic[921] <= 4'b0000;
        r_chickenpic[922] <= 4'b1111;
        r_chickenpic[923] <= 4'b1111;
        r_chickenpic[924] <= 4'b0000;
        r_chickenpic[925] <= 4'b0000;
        r_chickenpic[926] <= 4'b1111;
        r_chickenpic[927] <= 4'b1111;
        r_chickenpic[928] <= 4'b1111;
        r_chickenpic[929] <= 4'b1111;
        r_chickenpic[930] <= 4'b1111;
        r_chickenpic[931] <= 4'b1111;
        r_chickenpic[932] <= 4'b1111;
        r_chickenpic[933] <= 4'b1111;
        r_chickenpic[934] <= 4'b1111;
        r_chickenpic[935] <= 4'b1111;
        r_chickenpic[936] <= 4'b1111;
        r_chickenpic[937] <= 4'b1111;
        r_chickenpic[938] <= 4'b1111;
        r_chickenpic[939] <= 4'b1111;
        r_chickenpic[940] <= 4'b1111;
        r_chickenpic[941] <= 4'b1111;
        r_chickenpic[942] <= 4'b1111;
        r_chickenpic[943] <= 4'b1111;
        r_chickenpic[944] <= 4'b0000;
        r_chickenpic[945] <= 4'b0000;
        r_chickenpic[946] <= 4'b1111;
        r_chickenpic[947] <= 4'b1111;
        r_chickenpic[948] <= 4'b1111;
        r_chickenpic[949] <= 4'b1111;
        r_chickenpic[950] <= 4'b1111;
        r_chickenpic[951] <= 4'b1111;
        r_chickenpic[952] <= 4'b1111;
        r_chickenpic[953] <= 4'b1111;
        r_chickenpic[954] <= 4'b1111;
        r_chickenpic[955] <= 4'b1111;
        r_chickenpic[956] <= 4'b1111;
        r_chickenpic[957] <= 4'b1111;
        r_chickenpic[958] <= 4'b1111;
        r_chickenpic[959] <= 4'b1111;
        r_chickenpic[960] <= 4'b1111;
        r_chickenpic[961] <= 4'b1111;
        r_chickenpic[962] <= 4'b0000;
        r_chickenpic[963] <= 4'b0000;
        r_chickenpic[964] <= 4'b0000;
        r_chickenpic[965] <= 4'b0000;
        r_chickenpic[966] <= 4'b0000;
        r_chickenpic[967] <= 4'b0000;
        r_chickenpic[968] <= 4'b0000;
        r_chickenpic[969] <= 4'b0000;
        r_chickenpic[970] <= 4'b0000;
        r_chickenpic[971] <= 4'b0000;
        r_chickenpic[972] <= 4'b0000;
        r_chickenpic[973] <= 4'b0000;
        r_chickenpic[974] <= 4'b0000;
        r_chickenpic[975] <= 4'b1111;
        r_chickenpic[976] <= 4'b1111;
        r_chickenpic[977] <= 4'b1111;
        r_chickenpic[978] <= 4'b1111;
        r_chickenpic[979] <= 4'b1111;
        r_chickenpic[980] <= 4'b0000;
        r_chickenpic[981] <= 4'b0000;
        r_chickenpic[982] <= 4'b1111;
        r_chickenpic[983] <= 4'b1111;
        r_chickenpic[984] <= 4'b1111;
        r_chickenpic[985] <= 4'b1111;
        r_chickenpic[986] <= 4'b1111;
        r_chickenpic[987] <= 4'b1111;
        r_chickenpic[988] <= 4'b1111;
        r_chickenpic[989] <= 4'b1111;
        r_chickenpic[990] <= 4'b1111;
        r_chickenpic[991] <= 4'b1111;
        r_chickenpic[992] <= 4'b1111;
        r_chickenpic[993] <= 4'b1111;
        r_chickenpic[994] <= 4'b1111;
        r_chickenpic[995] <= 4'b1111;
        r_chickenpic[996] <= 4'b1111;
        r_chickenpic[997] <= 4'b1111;
        r_chickenpic[998] <= 4'b1111;
        r_chickenpic[999] <= 4'b0000;
        r_chickenpic[1000] <= 4'b1111;
        r_chickenpic[1001] <= 4'b1111;
        r_chickenpic[1002] <= 4'b1111;
        r_chickenpic[1003] <= 4'b1111;
        r_chickenpic[1004] <= 4'b1111;
        r_chickenpic[1005] <= 4'b1111;
        r_chickenpic[1006] <= 4'b1111;
        r_chickenpic[1007] <= 4'b1111;
        r_chickenpic[1008] <= 4'b1111;
        r_chickenpic[1009] <= 4'b1111;
        r_chickenpic[1010] <= 4'b1111;
        r_chickenpic[1011] <= 4'b1111;
        r_chickenpic[1012] <= 4'b1111;
        r_chickenpic[1013] <= 4'b1111;
        r_chickenpic[1014] <= 4'b1111;
        r_chickenpic[1015] <= 4'b1111;
        r_chickenpic[1016] <= 4'b1111;
        r_chickenpic[1017] <= 4'b0000;
        r_chickenpic[1018] <= 4'b0000;
        r_chickenpic[1019] <= 4'b0000;
        r_chickenpic[1020] <= 4'b0000;
        r_chickenpic[1021] <= 4'b0000;
        r_chickenpic[1022] <= 4'b0000;
        r_chickenpic[1023] <= 4'b0000;
        r_chickenpic[1024] <= 4'b0000;
        r_chickenpic[1025] <= 4'b0000;
        r_chickenpic[1026] <= 4'b0000;
        r_chickenpic[1027] <= 4'b0000;
        r_chickenpic[1028] <= 4'b1111;
        r_chickenpic[1029] <= 4'b1111;
        r_chickenpic[1030] <= 4'b1111;
        r_chickenpic[1031] <= 4'b1111;
        r_chickenpic[1032] <= 4'b1111;
        r_chickenpic[1033] <= 4'b1111;
        r_chickenpic[1034] <= 4'b1111;
        r_chickenpic[1035] <= 4'b0000;
        r_chickenpic[1036] <= 4'b0000;
        r_chickenpic[1037] <= 4'b1111;
        r_chickenpic[1038] <= 4'b1111;
        r_chickenpic[1039] <= 4'b1111;
        r_chickenpic[1040] <= 4'b1111;
        r_chickenpic[1041] <= 4'b1111;
        r_chickenpic[1042] <= 4'b1111;
        r_chickenpic[1043] <= 4'b1111;
        r_chickenpic[1044] <= 4'b1111;
        r_chickenpic[1045] <= 4'b1111;
        r_chickenpic[1046] <= 4'b1111;
        r_chickenpic[1047] <= 4'b1111;
        r_chickenpic[1048] <= 4'b1111;
        r_chickenpic[1049] <= 4'b1111;
        r_chickenpic[1050] <= 4'b1111;
        r_chickenpic[1051] <= 4'b1111;
        r_chickenpic[1052] <= 4'b1111;
        r_chickenpic[1053] <= 4'b0000;
        r_chickenpic[1054] <= 4'b0000;
        r_chickenpic[1055] <= 4'b1111;
        r_chickenpic[1056] <= 4'b1111;
        r_chickenpic[1057] <= 4'b1111;
        r_chickenpic[1058] <= 4'b1111;
        r_chickenpic[1059] <= 4'b1111;
        r_chickenpic[1060] <= 4'b1111;
        r_chickenpic[1061] <= 4'b1111;
        r_chickenpic[1062] <= 4'b1111;
        r_chickenpic[1063] <= 4'b1111;
        r_chickenpic[1064] <= 4'b1111;
        r_chickenpic[1065] <= 4'b1111;
        r_chickenpic[1066] <= 4'b1111;
        r_chickenpic[1067] <= 4'b1111;
        r_chickenpic[1068] <= 4'b1111;
        r_chickenpic[1069] <= 4'b1111;
        r_chickenpic[1070] <= 4'b1111;
        r_chickenpic[1071] <= 4'b1111;
        r_chickenpic[1072] <= 4'b0000;
        r_chickenpic[1073] <= 4'b0000;
        r_chickenpic[1074] <= 4'b1111;
        r_chickenpic[1075] <= 4'b1111;
        r_chickenpic[1076] <= 4'b1111;
        r_chickenpic[1077] <= 4'b1111;
        r_chickenpic[1078] <= 4'b1111;
        r_chickenpic[1079] <= 4'b1111;
        r_chickenpic[1080] <= 4'b1111;
        r_chickenpic[1081] <= 4'b1111;
        r_chickenpic[1082] <= 4'b1111;
        r_chickenpic[1083] <= 4'b1111;
        r_chickenpic[1084] <= 4'b1111;
        r_chickenpic[1085] <= 4'b1111;
        r_chickenpic[1086] <= 4'b1111;
        r_chickenpic[1087] <= 4'b1111;
        r_chickenpic[1088] <= 4'b1111;
        r_chickenpic[1089] <= 4'b1111;
        r_chickenpic[1090] <= 4'b0000;
        r_chickenpic[1091] <= 4'b0000;
        r_chickenpic[1092] <= 4'b1111;
        r_chickenpic[1093] <= 4'b1111;
        r_chickenpic[1094] <= 4'b1111;
        r_chickenpic[1095] <= 4'b1111;
        r_chickenpic[1096] <= 4'b1111;
        r_chickenpic[1097] <= 4'b1111;
        r_chickenpic[1098] <= 4'b1111;
        r_chickenpic[1099] <= 4'b1111;
        r_chickenpic[1100] <= 4'b1111;
        r_chickenpic[1101] <= 4'b1111;
        r_chickenpic[1102] <= 4'b1111;
        r_chickenpic[1103] <= 4'b1111;
        r_chickenpic[1104] <= 4'b1111;
        r_chickenpic[1105] <= 4'b1111;
        r_chickenpic[1106] <= 4'b1111;
        r_chickenpic[1107] <= 4'b1111;
        r_chickenpic[1108] <= 4'b0000;
        r_chickenpic[1109] <= 4'b0000;
        r_chickenpic[1110] <= 4'b1111;
        r_chickenpic[1111] <= 4'b1111;
        r_chickenpic[1112] <= 4'b1111;
        r_chickenpic[1113] <= 4'b1111;
        r_chickenpic[1114] <= 4'b1111;
        r_chickenpic[1115] <= 4'b1111;
        r_chickenpic[1116] <= 4'b1111;
        r_chickenpic[1117] <= 4'b1111;
        r_chickenpic[1118] <= 4'b1111;
        r_chickenpic[1119] <= 4'b1111;
        r_chickenpic[1120] <= 4'b1111;
        r_chickenpic[1121] <= 4'b1111;
        r_chickenpic[1122] <= 4'b1111;
        r_chickenpic[1123] <= 4'b1111;
        r_chickenpic[1124] <= 4'b1111;
        r_chickenpic[1125] <= 4'b1111;
        r_chickenpic[1126] <= 4'b1111;
        r_chickenpic[1127] <= 4'b0000;
        r_chickenpic[1128] <= 4'b0000;
        r_chickenpic[1129] <= 4'b1111;
        r_chickenpic[1130] <= 4'b1111;
        r_chickenpic[1131] <= 4'b1111;
        r_chickenpic[1132] <= 4'b1111;
        r_chickenpic[1133] <= 4'b1111;
        r_chickenpic[1134] <= 4'b1111;
        r_chickenpic[1135] <= 4'b1111;
        r_chickenpic[1136] <= 4'b1111;
        r_chickenpic[1137] <= 4'b1111;
        r_chickenpic[1138] <= 4'b1111;
        r_chickenpic[1139] <= 4'b1111;
        r_chickenpic[1140] <= 4'b1111;
        r_chickenpic[1141] <= 4'b1111;
        r_chickenpic[1142] <= 4'b1111;
        r_chickenpic[1143] <= 4'b1111;
        r_chickenpic[1144] <= 4'b1111;
        r_chickenpic[1145] <= 4'b1111;
        r_chickenpic[1146] <= 4'b0000;
        r_chickenpic[1147] <= 4'b1111;
        r_chickenpic[1148] <= 4'b1111;
        r_chickenpic[1149] <= 4'b1111;
        r_chickenpic[1150] <= 4'b1111;
        r_chickenpic[1151] <= 4'b1111;
        r_chickenpic[1152] <= 4'b1111;
        r_chickenpic[1153] <= 4'b1111;
        r_chickenpic[1154] <= 4'b1111;
        r_chickenpic[1155] <= 4'b1111;
        r_chickenpic[1156] <= 4'b1111;
        r_chickenpic[1157] <= 4'b1111;
        r_chickenpic[1158] <= 4'b1111;
        r_chickenpic[1159] <= 4'b1111;
        r_chickenpic[1160] <= 4'b1111;
        r_chickenpic[1161] <= 4'b1111;
        r_chickenpic[1162] <= 4'b1111;
        r_chickenpic[1163] <= 4'b0000;
        r_chickenpic[1164] <= 4'b0000;
        r_chickenpic[1165] <= 4'b1111;
        r_chickenpic[1166] <= 4'b1111;
        r_chickenpic[1167] <= 4'b1111;
        r_chickenpic[1168] <= 4'b1111;
        r_chickenpic[1169] <= 4'b1111;
        r_chickenpic[1170] <= 4'b1111;
        r_chickenpic[1171] <= 4'b1111;
        r_chickenpic[1172] <= 4'b1111;
        r_chickenpic[1173] <= 4'b1111;
        r_chickenpic[1174] <= 4'b1111;
        r_chickenpic[1175] <= 4'b1111;
        r_chickenpic[1176] <= 4'b1111;
        r_chickenpic[1177] <= 4'b1111;
        r_chickenpic[1178] <= 4'b1111;
        r_chickenpic[1179] <= 4'b1111;
        r_chickenpic[1180] <= 4'b1111;
        r_chickenpic[1181] <= 4'b1111;
        r_chickenpic[1182] <= 4'b0000;
        r_chickenpic[1183] <= 4'b1111;
        r_chickenpic[1184] <= 4'b1111;
        r_chickenpic[1185] <= 4'b1111;
        r_chickenpic[1186] <= 4'b1111;
        r_chickenpic[1187] <= 4'b1111;
        r_chickenpic[1188] <= 4'b1111;
        r_chickenpic[1189] <= 4'b1111;
        r_chickenpic[1190] <= 4'b1111;
        r_chickenpic[1191] <= 4'b1111;
        r_chickenpic[1192] <= 4'b1111;
        r_chickenpic[1193] <= 4'b1111;
        r_chickenpic[1194] <= 4'b1111;
        r_chickenpic[1195] <= 4'b1111;
        r_chickenpic[1196] <= 4'b1111;
        r_chickenpic[1197] <= 4'b1111;
        r_chickenpic[1198] <= 4'b1111;
        r_chickenpic[1199] <= 4'b1111;
        r_chickenpic[1200] <= 4'b1111;
        r_chickenpic[1201] <= 4'b0000;
        r_chickenpic[1202] <= 4'b1111;
        r_chickenpic[1203] <= 4'b1111;
        r_chickenpic[1204] <= 4'b1111;
        r_chickenpic[1205] <= 4'b1111;
        r_chickenpic[1206] <= 4'b1111;
        r_chickenpic[1207] <= 4'b1111;
        r_chickenpic[1208] <= 4'b1111;
        r_chickenpic[1209] <= 4'b1111;
        r_chickenpic[1210] <= 4'b1111;
        r_chickenpic[1211] <= 4'b1111;
        r_chickenpic[1212] <= 4'b1111;
        r_chickenpic[1213] <= 4'b1111;
        r_chickenpic[1214] <= 4'b1111;
        r_chickenpic[1215] <= 4'b1111;
        r_chickenpic[1216] <= 4'b1111;
        r_chickenpic[1217] <= 4'b1111;
        r_chickenpic[1218] <= 4'b0000;
        r_chickenpic[1219] <= 4'b1111;
        r_chickenpic[1220] <= 4'b1111;
        r_chickenpic[1221] <= 4'b1111;
        r_chickenpic[1222] <= 4'b1111;
        r_chickenpic[1223] <= 4'b1111;
        r_chickenpic[1224] <= 4'b1111;
        r_chickenpic[1225] <= 4'b1111;
        r_chickenpic[1226] <= 4'b1111;
        r_chickenpic[1227] <= 4'b1111;
        r_chickenpic[1228] <= 4'b1111;
        r_chickenpic[1229] <= 4'b1111;
        r_chickenpic[1230] <= 4'b1111;
        r_chickenpic[1231] <= 4'b1111;
        r_chickenpic[1232] <= 4'b1111;
        r_chickenpic[1233] <= 4'b1111;
        r_chickenpic[1234] <= 4'b1111;
        r_chickenpic[1235] <= 4'b1111;
        r_chickenpic[1236] <= 4'b0000;
        r_chickenpic[1237] <= 4'b0000;
        r_chickenpic[1238] <= 4'b1111;
        r_chickenpic[1239] <= 4'b1111;
        r_chickenpic[1240] <= 4'b1111;
        r_chickenpic[1241] <= 4'b1111;
        r_chickenpic[1242] <= 4'b1111;
        r_chickenpic[1243] <= 4'b1111;
        r_chickenpic[1244] <= 4'b1111;
        r_chickenpic[1245] <= 4'b1111;
        r_chickenpic[1246] <= 4'b1111;
        r_chickenpic[1247] <= 4'b1111;
        r_chickenpic[1248] <= 4'b1111;
        r_chickenpic[1249] <= 4'b1111;
        r_chickenpic[1250] <= 4'b1111;
        r_chickenpic[1251] <= 4'b1111;
        r_chickenpic[1252] <= 4'b1111;
        r_chickenpic[1253] <= 4'b1111;
        r_chickenpic[1254] <= 4'b1111;
        r_chickenpic[1255] <= 4'b1111;
        r_chickenpic[1256] <= 4'b0000;
        r_chickenpic[1257] <= 4'b1111;
        r_chickenpic[1258] <= 4'b1111;
        r_chickenpic[1259] <= 4'b1111;
        r_chickenpic[1260] <= 4'b1111;
        r_chickenpic[1261] <= 4'b1111;
        r_chickenpic[1262] <= 4'b1111;
        r_chickenpic[1263] <= 4'b1111;
        r_chickenpic[1264] <= 4'b1111;
        r_chickenpic[1265] <= 4'b1111;
        r_chickenpic[1266] <= 4'b1111;
        r_chickenpic[1267] <= 4'b1111;
        r_chickenpic[1268] <= 4'b1111;
        r_chickenpic[1269] <= 4'b1111;
        r_chickenpic[1270] <= 4'b1111;
        r_chickenpic[1271] <= 4'b1111;
        r_chickenpic[1272] <= 4'b1111;
        r_chickenpic[1273] <= 4'b0000;
        r_chickenpic[1274] <= 4'b1111;
        r_chickenpic[1275] <= 4'b1111;
        r_chickenpic[1276] <= 4'b1111;
        r_chickenpic[1277] <= 4'b1111;
        r_chickenpic[1278] <= 4'b1111;
        r_chickenpic[1279] <= 4'b1111;
        r_chickenpic[1280] <= 4'b1111;
        r_chickenpic[1281] <= 4'b1111;
        r_chickenpic[1282] <= 4'b1111;
        r_chickenpic[1283] <= 4'b1111;
        r_chickenpic[1284] <= 4'b1111;
        r_chickenpic[1285] <= 4'b1111;
        r_chickenpic[1286] <= 4'b1111;
        r_chickenpic[1287] <= 4'b1111;
        r_chickenpic[1288] <= 4'b1111;
        r_chickenpic[1289] <= 4'b1111;
        r_chickenpic[1290] <= 4'b1111;
        r_chickenpic[1291] <= 4'b0000;
        r_chickenpic[1292] <= 4'b0000;
        r_chickenpic[1293] <= 4'b1111;
        r_chickenpic[1294] <= 4'b1111;
        r_chickenpic[1295] <= 4'b1111;
        r_chickenpic[1296] <= 4'b1111;
        r_chickenpic[1297] <= 4'b0000;
        r_chickenpic[1298] <= 4'b1111;
        r_chickenpic[1299] <= 4'b1111;
        r_chickenpic[1300] <= 4'b1111;
        r_chickenpic[1301] <= 4'b1111;
        r_chickenpic[1302] <= 4'b1111;
        r_chickenpic[1303] <= 4'b1111;
        r_chickenpic[1304] <= 4'b1111;
        r_chickenpic[1305] <= 4'b1111;
        r_chickenpic[1306] <= 4'b1111;
        r_chickenpic[1307] <= 4'b1111;
        r_chickenpic[1308] <= 4'b1111;
        r_chickenpic[1309] <= 4'b1111;
        r_chickenpic[1310] <= 4'b1111;
        r_chickenpic[1311] <= 4'b0000;
        r_chickenpic[1312] <= 4'b1111;
        r_chickenpic[1313] <= 4'b1111;
        r_chickenpic[1314] <= 4'b1111;
        r_chickenpic[1315] <= 4'b1111;
        r_chickenpic[1316] <= 4'b1111;
        r_chickenpic[1317] <= 4'b1111;
        r_chickenpic[1318] <= 4'b1111;
        r_chickenpic[1319] <= 4'b1111;
        r_chickenpic[1320] <= 4'b1111;
        r_chickenpic[1321] <= 4'b1111;
        r_chickenpic[1322] <= 4'b1111;
        r_chickenpic[1323] <= 4'b1111;
        r_chickenpic[1324] <= 4'b1111;
        r_chickenpic[1325] <= 4'b1111;
        r_chickenpic[1326] <= 4'b1111;
        r_chickenpic[1327] <= 4'b1111;
        r_chickenpic[1328] <= 4'b0000;
        r_chickenpic[1329] <= 4'b1111;
        r_chickenpic[1330] <= 4'b1111;
        r_chickenpic[1331] <= 4'b1111;
        r_chickenpic[1332] <= 4'b1111;
        r_chickenpic[1333] <= 4'b1111;
        r_chickenpic[1334] <= 4'b1111;
        r_chickenpic[1335] <= 4'b1111;
        r_chickenpic[1336] <= 4'b1111;
        r_chickenpic[1337] <= 4'b1111;
        r_chickenpic[1338] <= 4'b1111;
        r_chickenpic[1339] <= 4'b1111;
        r_chickenpic[1340] <= 4'b1111;
        r_chickenpic[1341] <= 4'b1111;
        r_chickenpic[1342] <= 4'b1111;
        r_chickenpic[1343] <= 4'b1111;
        r_chickenpic[1344] <= 4'b1111;
        r_chickenpic[1345] <= 4'b0000;
        r_chickenpic[1346] <= 4'b0000;
        r_chickenpic[1347] <= 4'b1111;
        r_chickenpic[1348] <= 4'b1111;
        r_chickenpic[1349] <= 4'b1111;
        r_chickenpic[1350] <= 4'b1111;
        r_chickenpic[1351] <= 4'b0000;
        r_chickenpic[1352] <= 4'b0000;
        r_chickenpic[1353] <= 4'b0000;
        r_chickenpic[1354] <= 4'b0000;
        r_chickenpic[1355] <= 4'b1111;
        r_chickenpic[1356] <= 4'b1111;
        r_chickenpic[1357] <= 4'b1111;
        r_chickenpic[1358] <= 4'b1111;
        r_chickenpic[1359] <= 4'b1111;
        r_chickenpic[1360] <= 4'b1111;
        r_chickenpic[1361] <= 4'b1111;
        r_chickenpic[1362] <= 4'b1111;
        r_chickenpic[1363] <= 4'b1111;
        r_chickenpic[1364] <= 4'b1111;
        r_chickenpic[1365] <= 4'b1111;
        r_chickenpic[1366] <= 4'b0000;
        r_chickenpic[1367] <= 4'b1111;
        r_chickenpic[1368] <= 4'b1111;
        r_chickenpic[1369] <= 4'b1111;
        r_chickenpic[1370] <= 4'b1111;
        r_chickenpic[1371] <= 4'b1111;
        r_chickenpic[1372] <= 4'b1111;
        r_chickenpic[1373] <= 4'b1111;
        r_chickenpic[1374] <= 4'b1111;
        r_chickenpic[1375] <= 4'b1111;
        r_chickenpic[1376] <= 4'b1111;
        r_chickenpic[1377] <= 4'b1111;
        r_chickenpic[1378] <= 4'b1111;
        r_chickenpic[1379] <= 4'b1111;
        r_chickenpic[1380] <= 4'b1111;
        r_chickenpic[1381] <= 4'b1111;
        r_chickenpic[1382] <= 4'b1111;
        r_chickenpic[1383] <= 4'b0000;
        r_chickenpic[1384] <= 4'b1111;
        r_chickenpic[1385] <= 4'b1111;
        r_chickenpic[1386] <= 4'b1111;
        r_chickenpic[1387] <= 4'b1111;
        r_chickenpic[1388] <= 4'b1111;
        r_chickenpic[1389] <= 4'b1111;
        r_chickenpic[1390] <= 4'b1111;
        r_chickenpic[1391] <= 4'b1111;
        r_chickenpic[1392] <= 4'b1111;
        r_chickenpic[1393] <= 4'b1111;
        r_chickenpic[1394] <= 4'b1111;
        r_chickenpic[1395] <= 4'b1111;
        r_chickenpic[1396] <= 4'b1111;
        r_chickenpic[1397] <= 4'b1111;
        r_chickenpic[1398] <= 4'b1111;
        r_chickenpic[1399] <= 4'b0000;
        r_chickenpic[1400] <= 4'b0000;
        r_chickenpic[1401] <= 4'b1111;
        r_chickenpic[1402] <= 4'b1111;
        r_chickenpic[1403] <= 4'b1111;
        r_chickenpic[1404] <= 4'b1111;
        r_chickenpic[1405] <= 4'b1111;
        r_chickenpic[1406] <= 4'b1111;
        r_chickenpic[1407] <= 4'b1111;
        r_chickenpic[1408] <= 4'b1111;
        r_chickenpic[1409] <= 4'b0000;
        r_chickenpic[1410] <= 4'b0000;
        r_chickenpic[1411] <= 4'b0000;
        r_chickenpic[1412] <= 4'b1111;
        r_chickenpic[1413] <= 4'b1111;
        r_chickenpic[1414] <= 4'b1111;
        r_chickenpic[1415] <= 4'b1111;
        r_chickenpic[1416] <= 4'b1111;
        r_chickenpic[1417] <= 4'b1111;
        r_chickenpic[1418] <= 4'b1111;
        r_chickenpic[1419] <= 4'b1111;
        r_chickenpic[1420] <= 4'b0000;
        r_chickenpic[1421] <= 4'b0000;
        r_chickenpic[1422] <= 4'b1111;
        r_chickenpic[1423] <= 4'b1111;
        r_chickenpic[1424] <= 4'b1111;
        r_chickenpic[1425] <= 4'b1111;
        r_chickenpic[1426] <= 4'b1111;
        r_chickenpic[1427] <= 4'b1111;
        r_chickenpic[1428] <= 4'b1111;
        r_chickenpic[1429] <= 4'b1111;
        r_chickenpic[1430] <= 4'b1111;
        r_chickenpic[1431] <= 4'b1111;
        r_chickenpic[1432] <= 4'b1111;
        r_chickenpic[1433] <= 4'b1111;
        r_chickenpic[1434] <= 4'b1111;
        r_chickenpic[1435] <= 4'b1111;
        r_chickenpic[1436] <= 4'b1111;
        r_chickenpic[1437] <= 4'b1111;
        r_chickenpic[1438] <= 4'b0000;
        r_chickenpic[1439] <= 4'b1111;
        r_chickenpic[1440] <= 4'b1111;
        r_chickenpic[1441] <= 4'b1111;
        r_chickenpic[1442] <= 4'b1111;
        r_chickenpic[1443] <= 4'b1111;
        r_chickenpic[1444] <= 4'b1111;
        r_chickenpic[1445] <= 4'b1111;
        r_chickenpic[1446] <= 4'b1111;
        r_chickenpic[1447] <= 4'b1111;
        r_chickenpic[1448] <= 4'b1111;
        r_chickenpic[1449] <= 4'b1111;
        r_chickenpic[1450] <= 4'b1111;
        r_chickenpic[1451] <= 4'b1111;
        r_chickenpic[1452] <= 4'b1111;
        r_chickenpic[1453] <= 4'b0000;
        r_chickenpic[1454] <= 4'b0000;
        r_chickenpic[1455] <= 4'b1111;
        r_chickenpic[1456] <= 4'b1111;
        r_chickenpic[1457] <= 4'b1111;
        r_chickenpic[1458] <= 4'b1111;
        r_chickenpic[1459] <= 4'b1111;
        r_chickenpic[1460] <= 4'b1111;
        r_chickenpic[1461] <= 4'b1111;
        r_chickenpic[1462] <= 4'b1111;
        r_chickenpic[1463] <= 4'b1111;
        r_chickenpic[1464] <= 4'b1111;
        r_chickenpic[1465] <= 4'b0000;
        r_chickenpic[1466] <= 4'b0000;
        r_chickenpic[1467] <= 4'b0000;
        r_chickenpic[1468] <= 4'b1111;
        r_chickenpic[1469] <= 4'b1111;
        r_chickenpic[1470] <= 4'b1111;
        r_chickenpic[1471] <= 4'b1111;
        r_chickenpic[1472] <= 4'b1111;
        r_chickenpic[1473] <= 4'b1111;
        r_chickenpic[1474] <= 4'b1111;
        r_chickenpic[1475] <= 4'b0000;
        r_chickenpic[1476] <= 4'b0000;
        r_chickenpic[1477] <= 4'b1111;
        r_chickenpic[1478] <= 4'b1111;
        r_chickenpic[1479] <= 4'b1111;
        r_chickenpic[1480] <= 4'b1111;
        r_chickenpic[1481] <= 4'b1111;
        r_chickenpic[1482] <= 4'b1111;
        r_chickenpic[1483] <= 4'b1111;
        r_chickenpic[1484] <= 4'b1111;
        r_chickenpic[1485] <= 4'b1111;
        r_chickenpic[1486] <= 4'b1111;
        r_chickenpic[1487] <= 4'b1111;
        r_chickenpic[1488] <= 4'b1111;
        r_chickenpic[1489] <= 4'b1111;
        r_chickenpic[1490] <= 4'b1111;
        r_chickenpic[1491] <= 4'b1111;
        r_chickenpic[1492] <= 4'b1111;
        r_chickenpic[1493] <= 4'b0000;
        r_chickenpic[1494] <= 4'b0000;
        r_chickenpic[1495] <= 4'b1111;
        r_chickenpic[1496] <= 4'b1111;
        r_chickenpic[1497] <= 4'b1111;
        r_chickenpic[1498] <= 4'b1111;
        r_chickenpic[1499] <= 4'b1111;
        r_chickenpic[1500] <= 4'b1111;
        r_chickenpic[1501] <= 4'b1111;
        r_chickenpic[1502] <= 4'b1111;
        r_chickenpic[1503] <= 4'b1111;
        r_chickenpic[1504] <= 4'b1111;
        r_chickenpic[1505] <= 4'b1111;
        r_chickenpic[1506] <= 4'b1111;
        r_chickenpic[1507] <= 4'b0000;
        r_chickenpic[1508] <= 4'b0000;
        r_chickenpic[1509] <= 4'b1111;
        r_chickenpic[1510] <= 4'b1111;
        r_chickenpic[1511] <= 4'b1111;
        r_chickenpic[1512] <= 4'b1111;
        r_chickenpic[1513] <= 4'b1111;
        r_chickenpic[1514] <= 4'b1111;
        r_chickenpic[1515] <= 4'b1111;
        r_chickenpic[1516] <= 4'b1111;
        r_chickenpic[1517] <= 4'b1111;
        r_chickenpic[1518] <= 4'b1111;
        r_chickenpic[1519] <= 4'b1111;
        r_chickenpic[1520] <= 4'b0000;
        r_chickenpic[1521] <= 4'b0000;
        r_chickenpic[1522] <= 4'b0000;
        r_chickenpic[1523] <= 4'b0000;
        r_chickenpic[1524] <= 4'b1111;
        r_chickenpic[1525] <= 4'b1111;
        r_chickenpic[1526] <= 4'b1111;
        r_chickenpic[1527] <= 4'b1111;
        r_chickenpic[1528] <= 4'b1111;
        r_chickenpic[1529] <= 4'b1111;
        r_chickenpic[1530] <= 4'b0000;
        r_chickenpic[1531] <= 4'b0000;
        r_chickenpic[1532] <= 4'b1111;
        r_chickenpic[1533] <= 4'b1111;
        r_chickenpic[1534] <= 4'b1111;
        r_chickenpic[1535] <= 4'b1111;
        r_chickenpic[1536] <= 4'b1111;
        r_chickenpic[1537] <= 4'b1111;
        r_chickenpic[1538] <= 4'b1111;
        r_chickenpic[1539] <= 4'b1111;
        r_chickenpic[1540] <= 4'b1111;
        r_chickenpic[1541] <= 4'b1111;
        r_chickenpic[1542] <= 4'b1111;
        r_chickenpic[1543] <= 4'b1111;
        r_chickenpic[1544] <= 4'b1111;
        r_chickenpic[1545] <= 4'b1111;
        r_chickenpic[1546] <= 4'b1111;
        r_chickenpic[1547] <= 4'b1111;
        r_chickenpic[1548] <= 4'b0000;
        r_chickenpic[1549] <= 4'b0000;
        r_chickenpic[1550] <= 4'b1111;
        r_chickenpic[1551] <= 4'b1111;
        r_chickenpic[1552] <= 4'b1111;
        r_chickenpic[1553] <= 4'b1111;
        r_chickenpic[1554] <= 4'b1111;
        r_chickenpic[1555] <= 4'b1111;
        r_chickenpic[1556] <= 4'b1111;
        r_chickenpic[1557] <= 4'b1111;
        r_chickenpic[1558] <= 4'b1111;
        r_chickenpic[1559] <= 4'b1111;
        r_chickenpic[1560] <= 4'b1111;
        r_chickenpic[1561] <= 4'b1111;
        r_chickenpic[1562] <= 4'b1111;
        r_chickenpic[1563] <= 4'b1111;
        r_chickenpic[1564] <= 4'b1111;
        r_chickenpic[1565] <= 4'b1111;
        r_chickenpic[1566] <= 4'b1111;
        r_chickenpic[1567] <= 4'b1111;
        r_chickenpic[1568] <= 4'b1111;
        r_chickenpic[1569] <= 4'b1111;
        r_chickenpic[1570] <= 4'b1111;
        r_chickenpic[1571] <= 4'b1111;
        r_chickenpic[1572] <= 4'b1111;
        r_chickenpic[1573] <= 4'b0000;
        r_chickenpic[1574] <= 4'b0000;
        r_chickenpic[1575] <= 4'b0000;
        r_chickenpic[1576] <= 4'b1111;
        r_chickenpic[1577] <= 4'b1111;
        r_chickenpic[1578] <= 4'b0000;
        r_chickenpic[1579] <= 4'b0000;
        r_chickenpic[1580] <= 4'b1111;
        r_chickenpic[1581] <= 4'b1111;
        r_chickenpic[1582] <= 4'b1111;
        r_chickenpic[1583] <= 4'b1111;
        r_chickenpic[1584] <= 4'b1111;
        r_chickenpic[1585] <= 4'b0000;
        r_chickenpic[1586] <= 4'b0000;
        r_chickenpic[1587] <= 4'b1111;
        r_chickenpic[1588] <= 4'b1111;
        r_chickenpic[1589] <= 4'b1111;
        r_chickenpic[1590] <= 4'b1111;
        r_chickenpic[1591] <= 4'b1111;
        r_chickenpic[1592] <= 4'b1111;
        r_chickenpic[1593] <= 4'b1111;
        r_chickenpic[1594] <= 4'b1111;
        r_chickenpic[1595] <= 4'b1111;
        r_chickenpic[1596] <= 4'b1111;
        r_chickenpic[1597] <= 4'b1111;
        r_chickenpic[1598] <= 4'b1111;
        r_chickenpic[1599] <= 4'b1111;
        r_chickenpic[1600] <= 4'b1111;
        r_chickenpic[1601] <= 4'b1111;
        r_chickenpic[1602] <= 4'b1111;
        r_chickenpic[1603] <= 4'b0000;
        r_chickenpic[1604] <= 4'b0000;
        r_chickenpic[1605] <= 4'b1111;
        r_chickenpic[1606] <= 4'b1111;
        r_chickenpic[1607] <= 4'b1111;
        r_chickenpic[1608] <= 4'b1111;
        r_chickenpic[1609] <= 4'b1111;
        r_chickenpic[1610] <= 4'b1111;
        r_chickenpic[1611] <= 4'b1111;
        r_chickenpic[1612] <= 4'b1111;
        r_chickenpic[1613] <= 4'b1111;
        r_chickenpic[1614] <= 4'b1111;
        r_chickenpic[1615] <= 4'b1111;
        r_chickenpic[1616] <= 4'b1111;
        r_chickenpic[1617] <= 4'b1111;
        r_chickenpic[1618] <= 4'b1111;
        r_chickenpic[1619] <= 4'b1111;
        r_chickenpic[1620] <= 4'b1111;
        r_chickenpic[1621] <= 4'b1111;
        r_chickenpic[1622] <= 4'b1111;
        r_chickenpic[1623] <= 4'b1111;
        r_chickenpic[1624] <= 4'b1111;
        r_chickenpic[1625] <= 4'b1111;
        r_chickenpic[1626] <= 4'b1111;
        r_chickenpic[1627] <= 4'b1111;
        r_chickenpic[1628] <= 4'b1111;
        r_chickenpic[1629] <= 4'b0000;
        r_chickenpic[1630] <= 4'b0000;
        r_chickenpic[1631] <= 4'b0000;
        r_chickenpic[1632] <= 4'b0000;
        r_chickenpic[1633] <= 4'b1111;
        r_chickenpic[1634] <= 4'b0000;
        r_chickenpic[1635] <= 4'b1111;
        r_chickenpic[1636] <= 4'b1111;
        r_chickenpic[1637] <= 4'b1111;
        r_chickenpic[1638] <= 4'b1111;
        r_chickenpic[1639] <= 4'b1111;
        r_chickenpic[1640] <= 4'b0000;
        r_chickenpic[1641] <= 4'b1111;
        r_chickenpic[1642] <= 4'b1111;
        r_chickenpic[1643] <= 4'b1111;
        r_chickenpic[1644] <= 4'b1111;
        r_chickenpic[1645] <= 4'b1111;
        r_chickenpic[1646] <= 4'b1111;
        r_chickenpic[1647] <= 4'b1111;
        r_chickenpic[1648] <= 4'b1111;
        r_chickenpic[1649] <= 4'b1111;
        r_chickenpic[1650] <= 4'b1111;
        r_chickenpic[1651] <= 4'b1111;
        r_chickenpic[1652] <= 4'b1111;
        r_chickenpic[1653] <= 4'b1111;
        r_chickenpic[1654] <= 4'b1111;
        r_chickenpic[1655] <= 4'b1111;
        r_chickenpic[1656] <= 4'b1111;
        r_chickenpic[1657] <= 4'b1111;
        r_chickenpic[1658] <= 4'b1111;
        r_chickenpic[1659] <= 4'b0000;
        r_chickenpic[1660] <= 4'b1111;
        r_chickenpic[1661] <= 4'b1111;
        r_chickenpic[1662] <= 4'b1111;
        r_chickenpic[1663] <= 4'b1111;
        r_chickenpic[1664] <= 4'b1111;
        r_chickenpic[1665] <= 4'b1111;
        r_chickenpic[1666] <= 4'b1111;
        r_chickenpic[1667] <= 4'b1111;
        r_chickenpic[1668] <= 4'b1111;
        r_chickenpic[1669] <= 4'b1111;
        r_chickenpic[1670] <= 4'b1111;
        r_chickenpic[1671] <= 4'b1111;
        r_chickenpic[1672] <= 4'b1111;
        r_chickenpic[1673] <= 4'b1111;
        r_chickenpic[1674] <= 4'b1111;
        r_chickenpic[1675] <= 4'b1111;
        r_chickenpic[1676] <= 4'b1111;
        r_chickenpic[1677] <= 4'b1111;
        r_chickenpic[1678] <= 4'b1111;
        r_chickenpic[1679] <= 4'b1111;
        r_chickenpic[1680] <= 4'b1111;
        r_chickenpic[1681] <= 4'b1111;
        r_chickenpic[1682] <= 4'b0000;
        r_chickenpic[1683] <= 4'b0000;
        r_chickenpic[1684] <= 4'b0000;
        r_chickenpic[1685] <= 4'b1111;
        r_chickenpic[1686] <= 4'b1111;
        r_chickenpic[1687] <= 4'b0000;
        r_chickenpic[1688] <= 4'b0000;
        r_chickenpic[1689] <= 4'b0000;
        r_chickenpic[1690] <= 4'b0000;
        r_chickenpic[1691] <= 4'b1111;
        r_chickenpic[1692] <= 4'b1111;
        r_chickenpic[1693] <= 4'b1111;
        r_chickenpic[1694] <= 4'b0000;
        r_chickenpic[1695] <= 4'b0000;
        r_chickenpic[1696] <= 4'b1111;
        r_chickenpic[1697] <= 4'b1111;
        r_chickenpic[1698] <= 4'b1111;
        r_chickenpic[1699] <= 4'b1111;
        r_chickenpic[1700] <= 4'b1111;
        r_chickenpic[1701] <= 4'b1111;
        r_chickenpic[1702] <= 4'b1111;
        r_chickenpic[1703] <= 4'b1111;
        r_chickenpic[1704] <= 4'b1111;
        r_chickenpic[1705] <= 4'b1111;
        r_chickenpic[1706] <= 4'b1111;
        r_chickenpic[1707] <= 4'b1111;
        r_chickenpic[1708] <= 4'b1111;
        r_chickenpic[1709] <= 4'b1111;
        r_chickenpic[1710] <= 4'b1111;
        r_chickenpic[1711] <= 4'b1111;
        r_chickenpic[1712] <= 4'b1111;
        r_chickenpic[1713] <= 4'b1111;
        r_chickenpic[1714] <= 4'b0000;
        r_chickenpic[1715] <= 4'b0000;
        r_chickenpic[1716] <= 4'b1111;
        r_chickenpic[1717] <= 4'b1111;
        r_chickenpic[1718] <= 4'b1111;
        r_chickenpic[1719] <= 4'b1111;
        r_chickenpic[1720] <= 4'b1111;
        r_chickenpic[1721] <= 4'b1111;
        r_chickenpic[1722] <= 4'b1111;
        r_chickenpic[1723] <= 4'b1111;
        r_chickenpic[1724] <= 4'b1111;
        r_chickenpic[1725] <= 4'b1111;
        r_chickenpic[1726] <= 4'b1111;
        r_chickenpic[1727] <= 4'b1111;
        r_chickenpic[1728] <= 4'b1111;
        r_chickenpic[1729] <= 4'b1111;
        r_chickenpic[1730] <= 4'b1111;
        r_chickenpic[1731] <= 4'b1111;
        r_chickenpic[1732] <= 4'b1111;
        r_chickenpic[1733] <= 4'b1111;
        r_chickenpic[1734] <= 4'b1111;
        r_chickenpic[1735] <= 4'b1111;
        r_chickenpic[1736] <= 4'b1111;
        r_chickenpic[1737] <= 4'b0000;
        r_chickenpic[1738] <= 4'b0000;
        r_chickenpic[1739] <= 4'b0000;
        r_chickenpic[1740] <= 4'b1111;
        r_chickenpic[1741] <= 4'b1111;
        r_chickenpic[1742] <= 4'b1111;
        r_chickenpic[1743] <= 4'b0000;
        r_chickenpic[1744] <= 4'b0000;
        r_chickenpic[1745] <= 4'b0000;
        r_chickenpic[1746] <= 4'b1111;
        r_chickenpic[1747] <= 4'b1111;
        r_chickenpic[1748] <= 4'b1111;
        r_chickenpic[1749] <= 4'b0000;
        r_chickenpic[1750] <= 4'b0000;
        r_chickenpic[1751] <= 4'b1111;
        r_chickenpic[1752] <= 4'b1111;
        r_chickenpic[1753] <= 4'b1111;
        r_chickenpic[1754] <= 4'b1111;
        r_chickenpic[1755] <= 4'b1111;
        r_chickenpic[1756] <= 4'b1111;
        r_chickenpic[1757] <= 4'b1111;
        r_chickenpic[1758] <= 4'b1111;
        r_chickenpic[1759] <= 4'b1111;
        r_chickenpic[1760] <= 4'b1111;
        r_chickenpic[1761] <= 4'b1111;
        r_chickenpic[1762] <= 4'b1111;
        r_chickenpic[1763] <= 4'b1111;
        r_chickenpic[1764] <= 4'b1111;
        r_chickenpic[1765] <= 4'b1111;
        r_chickenpic[1766] <= 4'b1111;
        r_chickenpic[1767] <= 4'b1111;
        r_chickenpic[1768] <= 4'b1111;
        r_chickenpic[1769] <= 4'b1111;
        r_chickenpic[1770] <= 4'b0000;
        r_chickenpic[1771] <= 4'b1111;
        r_chickenpic[1772] <= 4'b1111;
        r_chickenpic[1773] <= 4'b1111;
        r_chickenpic[1774] <= 4'b1111;
        r_chickenpic[1775] <= 4'b1111;
        r_chickenpic[1776] <= 4'b1111;
        r_chickenpic[1777] <= 4'b1111;
        r_chickenpic[1778] <= 4'b1111;
        r_chickenpic[1779] <= 4'b1111;
        r_chickenpic[1780] <= 4'b1111;
        r_chickenpic[1781] <= 4'b1111;
        r_chickenpic[1782] <= 4'b1111;
        r_chickenpic[1783] <= 4'b1111;
        r_chickenpic[1784] <= 4'b1111;
        r_chickenpic[1785] <= 4'b1111;
        r_chickenpic[1786] <= 4'b1111;
        r_chickenpic[1787] <= 4'b1111;
        r_chickenpic[1788] <= 4'b1111;
        r_chickenpic[1789] <= 4'b1111;
        r_chickenpic[1790] <= 4'b1111;
        r_chickenpic[1791] <= 4'b1111;
        r_chickenpic[1792] <= 4'b0000;
        r_chickenpic[1793] <= 4'b1111;
        r_chickenpic[1794] <= 4'b1111;
        r_chickenpic[1795] <= 4'b0000;
        r_chickenpic[1796] <= 4'b0000;
        r_chickenpic[1797] <= 4'b0000;
        r_chickenpic[1798] <= 4'b0000;
        r_chickenpic[1799] <= 4'b0000;
        r_chickenpic[1800] <= 4'b0000;
        r_chickenpic[1801] <= 4'b1111;
        r_chickenpic[1802] <= 4'b1111;
        r_chickenpic[1803] <= 4'b0000;
        r_chickenpic[1804] <= 4'b0000;
        r_chickenpic[1805] <= 4'b1111;
        r_chickenpic[1806] <= 4'b1111;
        r_chickenpic[1807] <= 4'b1111;
        r_chickenpic[1808] <= 4'b1111;
        r_chickenpic[1809] <= 4'b1111;
        r_chickenpic[1810] <= 4'b1111;
        r_chickenpic[1811] <= 4'b1111;
        r_chickenpic[1812] <= 4'b1111;
        r_chickenpic[1813] <= 4'b1111;
        r_chickenpic[1814] <= 4'b1111;
        r_chickenpic[1815] <= 4'b1111;
        r_chickenpic[1816] <= 4'b1111;
        r_chickenpic[1817] <= 4'b1111;
        r_chickenpic[1818] <= 4'b1111;
        r_chickenpic[1819] <= 4'b1111;
        r_chickenpic[1820] <= 4'b1111;
        r_chickenpic[1821] <= 4'b1111;
        r_chickenpic[1822] <= 4'b1111;
        r_chickenpic[1823] <= 4'b1111;
        r_chickenpic[1824] <= 4'b1111;
        r_chickenpic[1825] <= 4'b0000;
        r_chickenpic[1826] <= 4'b0000;
        r_chickenpic[1827] <= 4'b1111;
        r_chickenpic[1828] <= 4'b1111;
        r_chickenpic[1829] <= 4'b1111;
        r_chickenpic[1830] <= 4'b1111;
        r_chickenpic[1831] <= 4'b1111;
        r_chickenpic[1832] <= 4'b1111;
        r_chickenpic[1833] <= 4'b1111;
        r_chickenpic[1834] <= 4'b1111;
        r_chickenpic[1835] <= 4'b1111;
        r_chickenpic[1836] <= 4'b1111;
        r_chickenpic[1837] <= 4'b1111;
        r_chickenpic[1838] <= 4'b1111;
        r_chickenpic[1839] <= 4'b1111;
        r_chickenpic[1840] <= 4'b1111;
        r_chickenpic[1841] <= 4'b1111;
        r_chickenpic[1842] <= 4'b1111;
        r_chickenpic[1843] <= 4'b1111;
        r_chickenpic[1844] <= 4'b0000;
        r_chickenpic[1845] <= 4'b0000;
        r_chickenpic[1846] <= 4'b0000;
        r_chickenpic[1847] <= 4'b0000;
        r_chickenpic[1848] <= 4'b1111;
        r_chickenpic[1849] <= 4'b1111;
        r_chickenpic[1850] <= 4'b1111;
        r_chickenpic[1851] <= 4'b1111;
        r_chickenpic[1852] <= 4'b1111;
        r_chickenpic[1853] <= 4'b0000;
        r_chickenpic[1854] <= 4'b0000;
        r_chickenpic[1855] <= 4'b0000;
        r_chickenpic[1856] <= 4'b1111;
        r_chickenpic[1857] <= 4'b1111;
        r_chickenpic[1858] <= 4'b0000;
        r_chickenpic[1859] <= 4'b0000;
        r_chickenpic[1860] <= 4'b1111;
        r_chickenpic[1861] <= 4'b1111;
        r_chickenpic[1862] <= 4'b1111;
        r_chickenpic[1863] <= 4'b1111;
        r_chickenpic[1864] <= 4'b1111;
        r_chickenpic[1865] <= 4'b1111;
        r_chickenpic[1866] <= 4'b1111;
        r_chickenpic[1867] <= 4'b1111;
        r_chickenpic[1868] <= 4'b1111;
        r_chickenpic[1869] <= 4'b1111;
        r_chickenpic[1870] <= 4'b1111;
        r_chickenpic[1871] <= 4'b1111;
        r_chickenpic[1872] <= 4'b1111;
        r_chickenpic[1873] <= 4'b1111;
        r_chickenpic[1874] <= 4'b1111;
        r_chickenpic[1875] <= 4'b1111;
        r_chickenpic[1876] <= 4'b1111;
        r_chickenpic[1877] <= 4'b1111;
        r_chickenpic[1878] <= 4'b1111;
        r_chickenpic[1879] <= 4'b1111;
        r_chickenpic[1880] <= 4'b1111;
        r_chickenpic[1881] <= 4'b0000;
        r_chickenpic[1882] <= 4'b0000;
        r_chickenpic[1883] <= 4'b1111;
        r_chickenpic[1884] <= 4'b1111;
        r_chickenpic[1885] <= 4'b1111;
        r_chickenpic[1886] <= 4'b1111;
        r_chickenpic[1887] <= 4'b1111;
        r_chickenpic[1888] <= 4'b1111;
        r_chickenpic[1889] <= 4'b1111;
        r_chickenpic[1890] <= 4'b1111;
        r_chickenpic[1891] <= 4'b1111;
        r_chickenpic[1892] <= 4'b1111;
        r_chickenpic[1893] <= 4'b1111;
        r_chickenpic[1894] <= 4'b0000;
        r_chickenpic[1895] <= 4'b0000;
        r_chickenpic[1896] <= 4'b1111;
        r_chickenpic[1897] <= 4'b1111;
        r_chickenpic[1898] <= 4'b1111;
        r_chickenpic[1899] <= 4'b0000;
        r_chickenpic[1900] <= 4'b0000;
        r_chickenpic[1901] <= 4'b0000;
        r_chickenpic[1902] <= 4'b0000;
        r_chickenpic[1903] <= 4'b0000;
        r_chickenpic[1904] <= 4'b0000;
        r_chickenpic[1905] <= 4'b0000;
        r_chickenpic[1906] <= 4'b0000;
        r_chickenpic[1907] <= 4'b0000;
        r_chickenpic[1908] <= 4'b0000;
        r_chickenpic[1909] <= 4'b0000;
        r_chickenpic[1910] <= 4'b1111;
        r_chickenpic[1911] <= 4'b1111;
        r_chickenpic[1912] <= 4'b0000;
        r_chickenpic[1913] <= 4'b0000;
        r_chickenpic[1914] <= 4'b1111;
        r_chickenpic[1915] <= 4'b1111;
        r_chickenpic[1916] <= 4'b1111;
        r_chickenpic[1917] <= 4'b1111;
        r_chickenpic[1918] <= 4'b1111;
        r_chickenpic[1919] <= 4'b1111;
        r_chickenpic[1920] <= 4'b1111;
        r_chickenpic[1921] <= 4'b1111;
        r_chickenpic[1922] <= 4'b1111;
        r_chickenpic[1923] <= 4'b1111;
        r_chickenpic[1924] <= 4'b1111;
        r_chickenpic[1925] <= 4'b1111;
        r_chickenpic[1926] <= 4'b1111;
        r_chickenpic[1927] <= 4'b1111;
        r_chickenpic[1928] <= 4'b1111;
        r_chickenpic[1929] <= 4'b1111;
        r_chickenpic[1930] <= 4'b1111;
        r_chickenpic[1931] <= 4'b1111;
        r_chickenpic[1932] <= 4'b1111;
        r_chickenpic[1933] <= 4'b1111;
        r_chickenpic[1934] <= 4'b1111;
        r_chickenpic[1935] <= 4'b1111;
        r_chickenpic[1936] <= 4'b1111;
        r_chickenpic[1937] <= 4'b0000;
        r_chickenpic[1938] <= 4'b0000;
        r_chickenpic[1939] <= 4'b1111;
        r_chickenpic[1940] <= 4'b1111;
        r_chickenpic[1941] <= 4'b1111;
        r_chickenpic[1942] <= 4'b1111;
        r_chickenpic[1943] <= 4'b1111;
        r_chickenpic[1944] <= 4'b1111;
        r_chickenpic[1945] <= 4'b1111;
        r_chickenpic[1946] <= 4'b1111;
        r_chickenpic[1947] <= 4'b1111;
        r_chickenpic[1948] <= 4'b1111;
        r_chickenpic[1949] <= 4'b1111;
        r_chickenpic[1950] <= 4'b0000;
        r_chickenpic[1951] <= 4'b0000;
        r_chickenpic[1952] <= 4'b0000;
        r_chickenpic[1953] <= 4'b1111;
        r_chickenpic[1954] <= 4'b0000;
        r_chickenpic[1955] <= 4'b0000;
        r_chickenpic[1956] <= 4'b1111;
        r_chickenpic[1957] <= 4'b1111;
        r_chickenpic[1958] <= 4'b1111;
        r_chickenpic[1959] <= 4'b0000;
        r_chickenpic[1960] <= 4'b0000;
        r_chickenpic[1961] <= 4'b0000;
        r_chickenpic[1962] <= 4'b0000;
        r_chickenpic[1963] <= 4'b0000;
        r_chickenpic[1964] <= 4'b1111;
        r_chickenpic[1965] <= 4'b1111;
        r_chickenpic[1966] <= 4'b0000;
        r_chickenpic[1967] <= 4'b0000;
        r_chickenpic[1968] <= 4'b1111;
        r_chickenpic[1969] <= 4'b1111;
        r_chickenpic[1970] <= 4'b1111;
        r_chickenpic[1971] <= 4'b1111;
        r_chickenpic[1972] <= 4'b1111;
        r_chickenpic[1973] <= 4'b1111;
        r_chickenpic[1974] <= 4'b1111;
        r_chickenpic[1975] <= 4'b1111;
        r_chickenpic[1976] <= 4'b1111;
        r_chickenpic[1977] <= 4'b1111;
        r_chickenpic[1978] <= 4'b1111;
        r_chickenpic[1979] <= 4'b1111;
        r_chickenpic[1980] <= 4'b1111;
        r_chickenpic[1981] <= 4'b1111;
        r_chickenpic[1982] <= 4'b1111;
        r_chickenpic[1983] <= 4'b1111;
        r_chickenpic[1984] <= 4'b1111;
        r_chickenpic[1985] <= 4'b1111;
        r_chickenpic[1986] <= 4'b1111;
        r_chickenpic[1987] <= 4'b1111;
        r_chickenpic[1988] <= 4'b1111;
        r_chickenpic[1989] <= 4'b1111;
        r_chickenpic[1990] <= 4'b1111;
        r_chickenpic[1991] <= 4'b1111;
        r_chickenpic[1992] <= 4'b0000;
        r_chickenpic[1993] <= 4'b0000;
        r_chickenpic[1994] <= 4'b0000;
        r_chickenpic[1995] <= 4'b1111;
        r_chickenpic[1996] <= 4'b1111;
        r_chickenpic[1997] <= 4'b1111;
        r_chickenpic[1998] <= 4'b1111;
        r_chickenpic[1999] <= 4'b1111;
        r_chickenpic[2000] <= 4'b1111;
        r_chickenpic[2001] <= 4'b1111;
        r_chickenpic[2002] <= 4'b1111;
        r_chickenpic[2003] <= 4'b1111;
        r_chickenpic[2004] <= 4'b1111;
        r_chickenpic[2005] <= 4'b1111;
        r_chickenpic[2006] <= 4'b0000;
        r_chickenpic[2007] <= 4'b0000;
        r_chickenpic[2008] <= 4'b0000;
        r_chickenpic[2009] <= 4'b0000;
        r_chickenpic[2010] <= 4'b0000;
        r_chickenpic[2011] <= 4'b0000;
        r_chickenpic[2012] <= 4'b0000;
        r_chickenpic[2013] <= 4'b0000;
        r_chickenpic[2014] <= 4'b0000;
        r_chickenpic[2015] <= 4'b0000;
        r_chickenpic[2016] <= 4'b1111;
        r_chickenpic[2017] <= 4'b1111;
        r_chickenpic[2018] <= 4'b1111;
        r_chickenpic[2019] <= 4'b1111;
        r_chickenpic[2020] <= 4'b1111;
        r_chickenpic[2021] <= 4'b0000;
        r_chickenpic[2022] <= 4'b0000;
        r_chickenpic[2023] <= 4'b1111;
        r_chickenpic[2024] <= 4'b1111;
        r_chickenpic[2025] <= 4'b1111;
        r_chickenpic[2026] <= 4'b1111;
        r_chickenpic[2027] <= 4'b1111;
        r_chickenpic[2028] <= 4'b1111;
        r_chickenpic[2029] <= 4'b1111;
        r_chickenpic[2030] <= 4'b1111;
        r_chickenpic[2031] <= 4'b1111;
        r_chickenpic[2032] <= 4'b1111;
        r_chickenpic[2033] <= 4'b1111;
        r_chickenpic[2034] <= 4'b1111;
        r_chickenpic[2035] <= 4'b1111;
        r_chickenpic[2036] <= 4'b1111;
        r_chickenpic[2037] <= 4'b1111;
        r_chickenpic[2038] <= 4'b1111;
        r_chickenpic[2039] <= 4'b1111;
        r_chickenpic[2040] <= 4'b1111;
        r_chickenpic[2041] <= 4'b1111;
        r_chickenpic[2042] <= 4'b1111;
        r_chickenpic[2043] <= 4'b1111;
        r_chickenpic[2044] <= 4'b1111;
        r_chickenpic[2045] <= 4'b1111;
        r_chickenpic[2046] <= 4'b1111;
        r_chickenpic[2047] <= 4'b1111;
        r_chickenpic[2048] <= 4'b0000;
        r_chickenpic[2049] <= 4'b0000;
        r_chickenpic[2050] <= 4'b0000;
        r_chickenpic[2051] <= 4'b1111;
        r_chickenpic[2052] <= 4'b1111;
        r_chickenpic[2053] <= 4'b1111;
        r_chickenpic[2054] <= 4'b1111;
        r_chickenpic[2055] <= 4'b1111;
        r_chickenpic[2056] <= 4'b1111;
        r_chickenpic[2057] <= 4'b1111;
        r_chickenpic[2058] <= 4'b1111;
        r_chickenpic[2059] <= 4'b1111;
        r_chickenpic[2060] <= 4'b1111;
        r_chickenpic[2061] <= 4'b1111;
        r_chickenpic[2062] <= 4'b1111;
        r_chickenpic[2063] <= 4'b1111;
        r_chickenpic[2064] <= 4'b0000;
        r_chickenpic[2065] <= 4'b0000;
        r_chickenpic[2066] <= 4'b0000;
        r_chickenpic[2067] <= 4'b1111;
        r_chickenpic[2068] <= 4'b1111;
        r_chickenpic[2069] <= 4'b1111;
        r_chickenpic[2070] <= 4'b1111;
        r_chickenpic[2071] <= 4'b1111;
        r_chickenpic[2072] <= 4'b1111;
        r_chickenpic[2073] <= 4'b1111;
        r_chickenpic[2074] <= 4'b1111;
        r_chickenpic[2075] <= 4'b0000;
        r_chickenpic[2076] <= 4'b0000;
        r_chickenpic[2077] <= 4'b1111;
        r_chickenpic[2078] <= 4'b1111;
        r_chickenpic[2079] <= 4'b1111;
        r_chickenpic[2080] <= 4'b1111;
        r_chickenpic[2081] <= 4'b1111;
        r_chickenpic[2082] <= 4'b1111;
        r_chickenpic[2083] <= 4'b1111;
        r_chickenpic[2084] <= 4'b1111;
        r_chickenpic[2085] <= 4'b1111;
        r_chickenpic[2086] <= 4'b1111;
        r_chickenpic[2087] <= 4'b1111;
        r_chickenpic[2088] <= 4'b1111;
        r_chickenpic[2089] <= 4'b1111;
        r_chickenpic[2090] <= 4'b1111;
        r_chickenpic[2091] <= 4'b1111;
        r_chickenpic[2092] <= 4'b1111;
        r_chickenpic[2093] <= 4'b1111;
        r_chickenpic[2094] <= 4'b1111;
        r_chickenpic[2095] <= 4'b1111;
        r_chickenpic[2096] <= 4'b1111;
        r_chickenpic[2097] <= 4'b1111;
        r_chickenpic[2098] <= 4'b1111;
        r_chickenpic[2099] <= 4'b1111;
        r_chickenpic[2100] <= 4'b1111;
        r_chickenpic[2101] <= 4'b1111;
        r_chickenpic[2102] <= 4'b1111;
        r_chickenpic[2103] <= 4'b1111;
        r_chickenpic[2104] <= 4'b0000;
        r_chickenpic[2105] <= 4'b0000;
        r_chickenpic[2106] <= 4'b0000;
        r_chickenpic[2107] <= 4'b1111;
        r_chickenpic[2108] <= 4'b1111;
        r_chickenpic[2109] <= 4'b1111;
        r_chickenpic[2110] <= 4'b1111;
        r_chickenpic[2111] <= 4'b1111;
        r_chickenpic[2112] <= 4'b1111;
        r_chickenpic[2113] <= 4'b1111;
        r_chickenpic[2114] <= 4'b1111;
        r_chickenpic[2115] <= 4'b1111;
        r_chickenpic[2116] <= 4'b1111;
        r_chickenpic[2117] <= 4'b1111;
        r_chickenpic[2118] <= 4'b1111;
        r_chickenpic[2119] <= 4'b1111;
        r_chickenpic[2120] <= 4'b1111;
        r_chickenpic[2121] <= 4'b1111;
        r_chickenpic[2122] <= 4'b1111;
        r_chickenpic[2123] <= 4'b1111;
        r_chickenpic[2124] <= 4'b1111;
        r_chickenpic[2125] <= 4'b1111;
        r_chickenpic[2126] <= 4'b1111;
        r_chickenpic[2127] <= 4'b1111;
        r_chickenpic[2128] <= 4'b0000;
        r_chickenpic[2129] <= 4'b0000;
        r_chickenpic[2130] <= 4'b0000;
        r_chickenpic[2131] <= 4'b1111;
        r_chickenpic[2132] <= 4'b1111;
        r_chickenpic[2133] <= 4'b1111;
        r_chickenpic[2134] <= 4'b1111;
        r_chickenpic[2135] <= 4'b1111;
        r_chickenpic[2136] <= 4'b1111;
        r_chickenpic[2137] <= 4'b1111;
        r_chickenpic[2138] <= 4'b1111;
        r_chickenpic[2139] <= 4'b1111;
        r_chickenpic[2140] <= 4'b1111;
        r_chickenpic[2141] <= 4'b1111;
        r_chickenpic[2142] <= 4'b1111;
        r_chickenpic[2143] <= 4'b1111;
        r_chickenpic[2144] <= 4'b1111;
        r_chickenpic[2145] <= 4'b1111;
        r_chickenpic[2146] <= 4'b1111;
        r_chickenpic[2147] <= 4'b1111;
        r_chickenpic[2148] <= 4'b1111;
        r_chickenpic[2149] <= 4'b1111;
        r_chickenpic[2150] <= 4'b1111;
        r_chickenpic[2151] <= 4'b1111;
        r_chickenpic[2152] <= 4'b1111;
        r_chickenpic[2153] <= 4'b1111;
        r_chickenpic[2154] <= 4'b1111;
        r_chickenpic[2155] <= 4'b1111;
        r_chickenpic[2156] <= 4'b1111;
        r_chickenpic[2157] <= 4'b1111;
        r_chickenpic[2158] <= 4'b1111;
        r_chickenpic[2159] <= 4'b1111;
        r_chickenpic[2160] <= 4'b1111;
        r_chickenpic[2161] <= 4'b0000;
        r_chickenpic[2162] <= 4'b0000;
        r_chickenpic[2163] <= 4'b0000;
        r_chickenpic[2164] <= 4'b1111;
        r_chickenpic[2165] <= 4'b1111;
        r_chickenpic[2166] <= 4'b1111;
        r_chickenpic[2167] <= 4'b1111;
        r_chickenpic[2168] <= 4'b1111;
        r_chickenpic[2169] <= 4'b1111;
        r_chickenpic[2170] <= 4'b1111;
        r_chickenpic[2171] <= 4'b1111;
        r_chickenpic[2172] <= 4'b1111;
        r_chickenpic[2173] <= 4'b1111;
        r_chickenpic[2174] <= 4'b1111;
        r_chickenpic[2175] <= 4'b1111;
        r_chickenpic[2176] <= 4'b1111;
        r_chickenpic[2177] <= 4'b1111;
        r_chickenpic[2178] <= 4'b1111;
        r_chickenpic[2179] <= 4'b1111;
        r_chickenpic[2180] <= 4'b1111;
        r_chickenpic[2181] <= 4'b1111;
        r_chickenpic[2182] <= 4'b0000;
        r_chickenpic[2183] <= 4'b0000;
        r_chickenpic[2184] <= 4'b0000;
        r_chickenpic[2185] <= 4'b1111;
        r_chickenpic[2186] <= 4'b1111;
        r_chickenpic[2187] <= 4'b1111;
        r_chickenpic[2188] <= 4'b1111;
        r_chickenpic[2189] <= 4'b1111;
        r_chickenpic[2190] <= 4'b1111;
        r_chickenpic[2191] <= 4'b1111;
        r_chickenpic[2192] <= 4'b1111;
        r_chickenpic[2193] <= 4'b1111;
        r_chickenpic[2194] <= 4'b1111;
        r_chickenpic[2195] <= 4'b1111;
        r_chickenpic[2196] <= 4'b1111;
        r_chickenpic[2197] <= 4'b1111;
        r_chickenpic[2198] <= 4'b1111;
        r_chickenpic[2199] <= 4'b1111;
        r_chickenpic[2200] <= 4'b1111;
        r_chickenpic[2201] <= 4'b1111;
        r_chickenpic[2202] <= 4'b1111;
        r_chickenpic[2203] <= 4'b1111;
        r_chickenpic[2204] <= 4'b1111;
        r_chickenpic[2205] <= 4'b1111;
        r_chickenpic[2206] <= 4'b1111;
        r_chickenpic[2207] <= 4'b1111;
        r_chickenpic[2208] <= 4'b1111;
        r_chickenpic[2209] <= 4'b1111;
        r_chickenpic[2210] <= 4'b1111;
        r_chickenpic[2211] <= 4'b1111;
        r_chickenpic[2212] <= 4'b1111;
        r_chickenpic[2213] <= 4'b1111;
        r_chickenpic[2214] <= 4'b1111;
        r_chickenpic[2215] <= 4'b1111;
        r_chickenpic[2216] <= 4'b1111;
        r_chickenpic[2217] <= 4'b0000;
        r_chickenpic[2218] <= 4'b0000;
        r_chickenpic[2219] <= 4'b0000;
        r_chickenpic[2220] <= 4'b0000;
        r_chickenpic[2221] <= 4'b1111;
        r_chickenpic[2222] <= 4'b1111;
        r_chickenpic[2223] <= 4'b1111;
        r_chickenpic[2224] <= 4'b1111;
        r_chickenpic[2225] <= 4'b1111;
        r_chickenpic[2226] <= 4'b1111;
        r_chickenpic[2227] <= 4'b1111;
        r_chickenpic[2228] <= 4'b1111;
        r_chickenpic[2229] <= 4'b1111;
        r_chickenpic[2230] <= 4'b1111;
        r_chickenpic[2231] <= 4'b1111;
        r_chickenpic[2232] <= 4'b1111;
        r_chickenpic[2233] <= 4'b1111;
        r_chickenpic[2234] <= 4'b0000;
        r_chickenpic[2235] <= 4'b0000;
        r_chickenpic[2236] <= 4'b0000;
        r_chickenpic[2237] <= 4'b0000;
        r_chickenpic[2238] <= 4'b0000;
        r_chickenpic[2239] <= 4'b1111;
        r_chickenpic[2240] <= 4'b1111;
        r_chickenpic[2241] <= 4'b1111;
        r_chickenpic[2242] <= 4'b1111;
        r_chickenpic[2243] <= 4'b1111;
        r_chickenpic[2244] <= 4'b1111;
        r_chickenpic[2245] <= 4'b1111;
        r_chickenpic[2246] <= 4'b1111;
        r_chickenpic[2247] <= 4'b1111;
        r_chickenpic[2248] <= 4'b1111;
        r_chickenpic[2249] <= 4'b1111;
        r_chickenpic[2250] <= 4'b1111;
        r_chickenpic[2251] <= 4'b1111;
        r_chickenpic[2252] <= 4'b1111;
        r_chickenpic[2253] <= 4'b1111;
        r_chickenpic[2254] <= 4'b1111;
        r_chickenpic[2255] <= 4'b1111;
        r_chickenpic[2256] <= 4'b1111;
        r_chickenpic[2257] <= 4'b1111;
        r_chickenpic[2258] <= 4'b1111;
        r_chickenpic[2259] <= 4'b1111;
        r_chickenpic[2260] <= 4'b1111;
        r_chickenpic[2261] <= 4'b1111;
        r_chickenpic[2262] <= 4'b1111;
        r_chickenpic[2263] <= 4'b1111;
        r_chickenpic[2264] <= 4'b1111;
        r_chickenpic[2265] <= 4'b1111;
        r_chickenpic[2266] <= 4'b1111;
        r_chickenpic[2267] <= 4'b1111;
        r_chickenpic[2268] <= 4'b1111;
        r_chickenpic[2269] <= 4'b1111;
        r_chickenpic[2270] <= 4'b1111;
        r_chickenpic[2271] <= 4'b1111;
        r_chickenpic[2272] <= 4'b1111;
        r_chickenpic[2273] <= 4'b1111;
        r_chickenpic[2274] <= 4'b0000;
        r_chickenpic[2275] <= 4'b0000;
        r_chickenpic[2276] <= 4'b0000;
        r_chickenpic[2277] <= 4'b0000;
        r_chickenpic[2278] <= 4'b0000;
        r_chickenpic[2279] <= 4'b0000;
        r_chickenpic[2280] <= 4'b1111;
        r_chickenpic[2281] <= 4'b1111;
        r_chickenpic[2282] <= 4'b1111;
        r_chickenpic[2283] <= 4'b1111;
        r_chickenpic[2284] <= 4'b1111;
        r_chickenpic[2285] <= 4'b1111;
        r_chickenpic[2286] <= 4'b0000;
        r_chickenpic[2287] <= 4'b0000;
        r_chickenpic[2288] <= 4'b0000;
        r_chickenpic[2289] <= 4'b0000;
        r_chickenpic[2290] <= 4'b0000;
        r_chickenpic[2291] <= 4'b0000;
        r_chickenpic[2292] <= 4'b0000;
        r_chickenpic[2293] <= 4'b1111;
        r_chickenpic[2294] <= 4'b1111;
        r_chickenpic[2295] <= 4'b1111;
        r_chickenpic[2296] <= 4'b1111;
        r_chickenpic[2297] <= 4'b1111;
        r_chickenpic[2298] <= 4'b1111;
        r_chickenpic[2299] <= 4'b1111;
        r_chickenpic[2300] <= 4'b1111;
        r_chickenpic[2301] <= 4'b1111;
        r_chickenpic[2302] <= 4'b1111;
        r_chickenpic[2303] <= 4'b1111;
        r_chickenpic[2304] <= 4'b1111;
        r_chickenpic[2305] <= 4'b1111;
        r_chickenpic[2306] <= 4'b1111;
        r_chickenpic[2307] <= 4'b1111;
        r_chickenpic[2308] <= 4'b1111;
        r_chickenpic[2309] <= 4'b1111;
        r_chickenpic[2310] <= 4'b1111;
        r_chickenpic[2311] <= 4'b1111;
        r_chickenpic[2312] <= 4'b1111;
        r_chickenpic[2313] <= 4'b1111;
        r_chickenpic[2314] <= 4'b1111;
        r_chickenpic[2315] <= 4'b1111;
        r_chickenpic[2316] <= 4'b1111;
        r_chickenpic[2317] <= 4'b1111;
        r_chickenpic[2318] <= 4'b1111;
        r_chickenpic[2319] <= 4'b1111;
        r_chickenpic[2320] <= 4'b1111;
        r_chickenpic[2321] <= 4'b1111;
        r_chickenpic[2322] <= 4'b1111;
        r_chickenpic[2323] <= 4'b1111;
        r_chickenpic[2324] <= 4'b1111;
        r_chickenpic[2325] <= 4'b1111;
        r_chickenpic[2326] <= 4'b1111;
        r_chickenpic[2327] <= 4'b1111;
        r_chickenpic[2328] <= 4'b1111;
        r_chickenpic[2329] <= 4'b1111;
        r_chickenpic[2330] <= 4'b0000;
        r_chickenpic[2331] <= 4'b0000;
        r_chickenpic[2332] <= 4'b0000;
        r_chickenpic[2333] <= 4'b0000;
        r_chickenpic[2334] <= 4'b0000;
        r_chickenpic[2335] <= 4'b0000;
        r_chickenpic[2336] <= 4'b0000;
        r_chickenpic[2337] <= 4'b0000;
        r_chickenpic[2338] <= 4'b0000;
        r_chickenpic[2339] <= 4'b0000;
        r_chickenpic[2340] <= 4'b0000;
        r_chickenpic[2341] <= 4'b0000;
        r_chickenpic[2342] <= 4'b0000;
        r_chickenpic[2343] <= 4'b0000;
        r_chickenpic[2344] <= 4'b0000;
        r_chickenpic[2345] <= 4'b1111;
        r_chickenpic[2346] <= 4'b0000;
        r_chickenpic[2347] <= 4'b1111;
        r_chickenpic[2348] <= 4'b1111;
        r_chickenpic[2349] <= 4'b1111;
        r_chickenpic[2350] <= 4'b1111;
        r_chickenpic[2351] <= 4'b1111;
        r_chickenpic[2352] <= 4'b1111;
        r_chickenpic[2353] <= 4'b1111;
        r_chickenpic[2354] <= 4'b1111;
        r_chickenpic[2355] <= 4'b1111;
        r_chickenpic[2356] <= 4'b1111;
        r_chickenpic[2357] <= 4'b1111;
        r_chickenpic[2358] <= 4'b1111;
        r_chickenpic[2359] <= 4'b1111;
        r_chickenpic[2360] <= 4'b1111;
        r_chickenpic[2361] <= 4'b1111;
        r_chickenpic[2362] <= 4'b1111;
        r_chickenpic[2363] <= 4'b1111;
        r_chickenpic[2364] <= 4'b1111;
        r_chickenpic[2365] <= 4'b1111;
        r_chickenpic[2366] <= 4'b1111;
        r_chickenpic[2367] <= 4'b1111;
        r_chickenpic[2368] <= 4'b1111;
        r_chickenpic[2369] <= 4'b1111;
        r_chickenpic[2370] <= 4'b1111;
        r_chickenpic[2371] <= 4'b1111;
        r_chickenpic[2372] <= 4'b1111;
        r_chickenpic[2373] <= 4'b1111;
        r_chickenpic[2374] <= 4'b1111;
        r_chickenpic[2375] <= 4'b1111;
        r_chickenpic[2376] <= 4'b1111;
        r_chickenpic[2377] <= 4'b1111;
        r_chickenpic[2378] <= 4'b1111;
        r_chickenpic[2379] <= 4'b1111;
        r_chickenpic[2380] <= 4'b1111;
        r_chickenpic[2381] <= 4'b1111;
        r_chickenpic[2382] <= 4'b1111;
        r_chickenpic[2383] <= 4'b1111;
        r_chickenpic[2384] <= 4'b1111;
        r_chickenpic[2385] <= 4'b0000;
        r_chickenpic[2386] <= 4'b0000;
        r_chickenpic[2387] <= 4'b0000;
        r_chickenpic[2388] <= 4'b1111;
        r_chickenpic[2389] <= 4'b1111;
        r_chickenpic[2390] <= 4'b1111;
        r_chickenpic[2391] <= 4'b1111;
        r_chickenpic[2392] <= 4'b1111;
        r_chickenpic[2393] <= 4'b1111;
        r_chickenpic[2394] <= 4'b1111;
        r_chickenpic[2395] <= 4'b1111;
        r_chickenpic[2396] <= 4'b1111;
        r_chickenpic[2397] <= 4'b1111;
        r_chickenpic[2398] <= 4'b0000;
        r_chickenpic[2399] <= 4'b0000;
        r_chickenpic[2400] <= 4'b0000;
        r_chickenpic[2401] <= 4'b0000;
        r_chickenpic[2402] <= 4'b1111;
        r_chickenpic[2403] <= 4'b1111;
        r_chickenpic[2404] <= 4'b1111;
        r_chickenpic[2405] <= 4'b1111;
        r_chickenpic[2406] <= 4'b1111;
        r_chickenpic[2407] <= 4'b1111;
        r_chickenpic[2408] <= 4'b1111;
        r_chickenpic[2409] <= 4'b1111;
        r_chickenpic[2410] <= 4'b1111;
        r_chickenpic[2411] <= 4'b1111;
        r_chickenpic[2412] <= 4'b1111;
        r_chickenpic[2413] <= 4'b1111;
        r_chickenpic[2414] <= 4'b1111;
        r_chickenpic[2415] <= 4'b1111;
        r_chickenpic[2416] <= 4'b1111;
        r_chickenpic[2417] <= 4'b1111;
        r_chickenpic[2418] <= 4'b1111;
        r_chickenpic[2419] <= 4'b1111;
        r_chickenpic[2420] <= 4'b1111;
        r_chickenpic[2421] <= 4'b1111;
        r_chickenpic[2422] <= 4'b1111;
        r_chickenpic[2423] <= 4'b1111;
        r_chickenpic[2424] <= 4'b1111;
        r_chickenpic[2425] <= 4'b1111;
        r_chickenpic[2426] <= 4'b1111;
        r_chickenpic[2427] <= 4'b1111;
        r_chickenpic[2428] <= 4'b1111;
        r_chickenpic[2429] <= 4'b1111;
        r_chickenpic[2430] <= 4'b1111;
        r_chickenpic[2431] <= 4'b1111;
        r_chickenpic[2432] <= 4'b1111;
        r_chickenpic[2433] <= 4'b1111;
        r_chickenpic[2434] <= 4'b0000;
        r_chickenpic[2435] <= 4'b1111;
        r_chickenpic[2436] <= 4'b1111;
        r_chickenpic[2437] <= 4'b1111;
        r_chickenpic[2438] <= 4'b1111;
        r_chickenpic[2439] <= 4'b1111;
        r_chickenpic[2440] <= 4'b0000;
        r_chickenpic[2441] <= 4'b0000;
        r_chickenpic[2442] <= 4'b1111;
        r_chickenpic[2443] <= 4'b1111;
        r_chickenpic[2444] <= 4'b1111;
        r_chickenpic[2445] <= 4'b1111;
        r_chickenpic[2446] <= 4'b1111;
        r_chickenpic[2447] <= 4'b1111;
        r_chickenpic[2448] <= 4'b1111;
        r_chickenpic[2449] <= 4'b1111;
        r_chickenpic[2450] <= 4'b1111;
        r_chickenpic[2451] <= 4'b1111;
        r_chickenpic[2452] <= 4'b1111;
        r_chickenpic[2453] <= 4'b0000;
        r_chickenpic[2454] <= 4'b0000;
        r_chickenpic[2455] <= 4'b0000;
        r_chickenpic[2456] <= 4'b1111;
        r_chickenpic[2457] <= 4'b1111;
        r_chickenpic[2458] <= 4'b1111;
        r_chickenpic[2459] <= 4'b1111;
        r_chickenpic[2460] <= 4'b1111;
        r_chickenpic[2461] <= 4'b1111;
        r_chickenpic[2462] <= 4'b1111;
        r_chickenpic[2463] <= 4'b1111;
        r_chickenpic[2464] <= 4'b1111;
        r_chickenpic[2465] <= 4'b1111;
        r_chickenpic[2466] <= 4'b1111;
        r_chickenpic[2467] <= 4'b1111;
        r_chickenpic[2468] <= 4'b1111;
        r_chickenpic[2469] <= 4'b1111;
        r_chickenpic[2470] <= 4'b1111;
        r_chickenpic[2471] <= 4'b1111;
        r_chickenpic[2472] <= 4'b1111;
        r_chickenpic[2473] <= 4'b1111;
        r_chickenpic[2474] <= 4'b1111;
        r_chickenpic[2475] <= 4'b1111;
        r_chickenpic[2476] <= 4'b1111;
        r_chickenpic[2477] <= 4'b1111;
        r_chickenpic[2478] <= 4'b1111;
        r_chickenpic[2479] <= 4'b1111;
        r_chickenpic[2480] <= 4'b1111;
        r_chickenpic[2481] <= 4'b1111;
        r_chickenpic[2482] <= 4'b1111;
        r_chickenpic[2483] <= 4'b1111;
        r_chickenpic[2484] <= 4'b1111;
        r_chickenpic[2485] <= 4'b1111;
        r_chickenpic[2486] <= 4'b1111;
        r_chickenpic[2487] <= 4'b1111;
        r_chickenpic[2488] <= 4'b1111;
        r_chickenpic[2489] <= 4'b0000;
        r_chickenpic[2490] <= 4'b0000;
        r_chickenpic[2491] <= 4'b0000;
        r_chickenpic[2492] <= 4'b0000;
        r_chickenpic[2493] <= 4'b0000;
        r_chickenpic[2494] <= 4'b0000;
        r_chickenpic[2495] <= 4'b0000;
        r_chickenpic[2496] <= 4'b0000;
        r_chickenpic[2497] <= 4'b0000;
        r_chickenpic[2498] <= 4'b0000;
        r_chickenpic[2499] <= 4'b0000;
        r_chickenpic[2500] <= 4'b1111;
        r_chickenpic[2501] <= 4'b1111;
        r_chickenpic[2502] <= 4'b0000;
        r_chickenpic[2503] <= 4'b0000;
        r_chickenpic[2504] <= 4'b1111;
        r_chickenpic[2505] <= 4'b1111;
        r_chickenpic[2506] <= 4'b1111;
        r_chickenpic[2507] <= 4'b0000;
        r_chickenpic[2508] <= 4'b0000;
        r_chickenpic[2509] <= 4'b0000;
        r_chickenpic[2510] <= 4'b0000;
        r_chickenpic[2511] <= 4'b1111;
        r_chickenpic[2512] <= 4'b1111;
        r_chickenpic[2513] <= 4'b0000;
        r_chickenpic[2514] <= 4'b1111;
        r_chickenpic[2515] <= 4'b1111;
        r_chickenpic[2516] <= 4'b1111;
        r_chickenpic[2517] <= 4'b1111;
        r_chickenpic[2518] <= 4'b1111;
        r_chickenpic[2519] <= 4'b1111;
        r_chickenpic[2520] <= 4'b1111;
        r_chickenpic[2521] <= 4'b1111;
        r_chickenpic[2522] <= 4'b1111;
        r_chickenpic[2523] <= 4'b1111;
        r_chickenpic[2524] <= 4'b1111;
        r_chickenpic[2525] <= 4'b1111;
        r_chickenpic[2526] <= 4'b1111;
        r_chickenpic[2527] <= 4'b1111;
        r_chickenpic[2528] <= 4'b1111;
        r_chickenpic[2529] <= 4'b1111;
        r_chickenpic[2530] <= 4'b1111;
        r_chickenpic[2531] <= 4'b1111;
        r_chickenpic[2532] <= 4'b1111;
        r_chickenpic[2533] <= 4'b1111;
        r_chickenpic[2534] <= 4'b1111;
        r_chickenpic[2535] <= 4'b1111;
        r_chickenpic[2536] <= 4'b1111;
        r_chickenpic[2537] <= 4'b1111;
        r_chickenpic[2538] <= 4'b1111;
        r_chickenpic[2539] <= 4'b1111;
        r_chickenpic[2540] <= 4'b1111;
        r_chickenpic[2541] <= 4'b1111;
        r_chickenpic[2542] <= 4'b1111;
        r_chickenpic[2543] <= 4'b0000;
        r_chickenpic[2544] <= 4'b0000;
        r_chickenpic[2545] <= 4'b0000;
        r_chickenpic[2546] <= 4'b0000;
        r_chickenpic[2547] <= 4'b0000;
        r_chickenpic[2548] <= 4'b0000;
        r_chickenpic[2549] <= 4'b0000;
        r_chickenpic[2550] <= 4'b1111;
        r_chickenpic[2551] <= 4'b0000;
        r_chickenpic[2552] <= 4'b0000;
        r_chickenpic[2553] <= 4'b1111;
        r_chickenpic[2554] <= 4'b1111;
        r_chickenpic[2555] <= 4'b1111;
        r_chickenpic[2556] <= 4'b1111;
        r_chickenpic[2557] <= 4'b1111;
        r_chickenpic[2558] <= 4'b0000;
        r_chickenpic[2559] <= 4'b0000;
        r_chickenpic[2560] <= 4'b0000;
        r_chickenpic[2561] <= 4'b0000;
        r_chickenpic[2562] <= 4'b0000;
        r_chickenpic[2563] <= 4'b0000;
        r_chickenpic[2564] <= 4'b0000;
        r_chickenpic[2565] <= 4'b0000;
        r_chickenpic[2566] <= 4'b0000;
        r_chickenpic[2567] <= 4'b0000;
        r_chickenpic[2568] <= 4'b1111;
        r_chickenpic[2569] <= 4'b1111;
        r_chickenpic[2570] <= 4'b1111;
        r_chickenpic[2571] <= 4'b1111;
        r_chickenpic[2572] <= 4'b1111;
        r_chickenpic[2573] <= 4'b1111;
        r_chickenpic[2574] <= 4'b1111;
        r_chickenpic[2575] <= 4'b1111;
        r_chickenpic[2576] <= 4'b1111;
        r_chickenpic[2577] <= 4'b1111;
        r_chickenpic[2578] <= 4'b1111;
        r_chickenpic[2579] <= 4'b1111;
        r_chickenpic[2580] <= 4'b1111;
        r_chickenpic[2581] <= 4'b1111;
        r_chickenpic[2582] <= 4'b1111;
        r_chickenpic[2583] <= 4'b1111;
        r_chickenpic[2584] <= 4'b1111;
        r_chickenpic[2585] <= 4'b1111;
        r_chickenpic[2586] <= 4'b1111;
        r_chickenpic[2587] <= 4'b1111;
        r_chickenpic[2588] <= 4'b1111;
        r_chickenpic[2589] <= 4'b1111;
        r_chickenpic[2590] <= 4'b1111;
        r_chickenpic[2591] <= 4'b1111;
        r_chickenpic[2592] <= 4'b1111;
        r_chickenpic[2593] <= 4'b1111;
        r_chickenpic[2594] <= 4'b1111;
        r_chickenpic[2595] <= 4'b1111;
        r_chickenpic[2596] <= 4'b1111;
        r_chickenpic[2597] <= 4'b1111;
        r_chickenpic[2598] <= 4'b1111;
        r_chickenpic[2599] <= 4'b0000;
        r_chickenpic[2600] <= 4'b0000;
        r_chickenpic[2601] <= 4'b0000;
        r_chickenpic[2602] <= 4'b0000;
        r_chickenpic[2603] <= 4'b0000;
        r_chickenpic[2604] <= 4'b1111;
        r_chickenpic[2605] <= 4'b1111;
        r_chickenpic[2606] <= 4'b1111;
        r_chickenpic[2607] <= 4'b1111;
        r_chickenpic[2608] <= 4'b1111;
        r_chickenpic[2609] <= 4'b1111;
        r_chickenpic[2610] <= 4'b1111;
        r_chickenpic[2611] <= 4'b1111;
        r_chickenpic[2612] <= 4'b0000;
        r_chickenpic[2613] <= 4'b0000;
        r_chickenpic[2614] <= 4'b0000;
        r_chickenpic[2615] <= 4'b0000;
        r_chickenpic[2616] <= 4'b0000;
        r_chickenpic[2617] <= 4'b0000;
        r_chickenpic[2618] <= 4'b1111;
        r_chickenpic[2619] <= 4'b1111;
        r_chickenpic[2620] <= 4'b1111;
        r_chickenpic[2621] <= 4'b0000;
        r_chickenpic[2622] <= 4'b1111;
        r_chickenpic[2623] <= 4'b1111;
        r_chickenpic[2624] <= 4'b1111;
        r_chickenpic[2625] <= 4'b1111;
        r_chickenpic[2626] <= 4'b1111;
        r_chickenpic[2627] <= 4'b1111;
        r_chickenpic[2628] <= 4'b1111;
        r_chickenpic[2629] <= 4'b1111;
        r_chickenpic[2630] <= 4'b1111;
        r_chickenpic[2631] <= 4'b1111;
        r_chickenpic[2632] <= 4'b1111;
        r_chickenpic[2633] <= 4'b1111;
        r_chickenpic[2634] <= 4'b1111;
        r_chickenpic[2635] <= 4'b1111;
        r_chickenpic[2636] <= 4'b1111;
        r_chickenpic[2637] <= 4'b1111;
        r_chickenpic[2638] <= 4'b1111;
        r_chickenpic[2639] <= 4'b1111;
        r_chickenpic[2640] <= 4'b1111;
        r_chickenpic[2641] <= 4'b1111;
        r_chickenpic[2642] <= 4'b1111;
        r_chickenpic[2643] <= 4'b1111;
        r_chickenpic[2644] <= 4'b1111;
        r_chickenpic[2645] <= 4'b1111;
        r_chickenpic[2646] <= 4'b1111;
        r_chickenpic[2647] <= 4'b1111;
        r_chickenpic[2648] <= 4'b1111;
        r_chickenpic[2649] <= 4'b1111;
        r_chickenpic[2650] <= 4'b1111;
        r_chickenpic[2651] <= 4'b1111;
        r_chickenpic[2652] <= 4'b1111;
        r_chickenpic[2653] <= 4'b1111;
        r_chickenpic[2654] <= 4'b0000;
        r_chickenpic[2655] <= 4'b0000;
        r_chickenpic[2656] <= 4'b0000;
        r_chickenpic[2657] <= 4'b0000;
        r_chickenpic[2658] <= 4'b1111;
        r_chickenpic[2659] <= 4'b1111;
        r_chickenpic[2660] <= 4'b1111;
        r_chickenpic[2661] <= 4'b1111;
        r_chickenpic[2662] <= 4'b1111;
        r_chickenpic[2663] <= 4'b1111;
        r_chickenpic[2664] <= 4'b1111;
        r_chickenpic[2665] <= 4'b1111;
        r_chickenpic[2666] <= 4'b1111;
        r_chickenpic[2667] <= 4'b0000;
        r_chickenpic[2668] <= 4'b0000;
        r_chickenpic[2669] <= 4'b0000;
        r_chickenpic[2670] <= 4'b0000;
        r_chickenpic[2671] <= 4'b0000;
        r_chickenpic[2672] <= 4'b1111;
        r_chickenpic[2673] <= 4'b1111;
        r_chickenpic[2674] <= 4'b1111;
        r_chickenpic[2675] <= 4'b1111;
        r_chickenpic[2676] <= 4'b1111;
        r_chickenpic[2677] <= 4'b1111;
        r_chickenpic[2678] <= 4'b1111;
        r_chickenpic[2679] <= 4'b1111;
        r_chickenpic[2680] <= 4'b1111;
        r_chickenpic[2681] <= 4'b1111;
        r_chickenpic[2682] <= 4'b1111;
        r_chickenpic[2683] <= 4'b1111;
        r_chickenpic[2684] <= 4'b1111;
        r_chickenpic[2685] <= 4'b1111;
        r_chickenpic[2686] <= 4'b1111;
        r_chickenpic[2687] <= 4'b1111;
        r_chickenpic[2688] <= 4'b1111;
        r_chickenpic[2689] <= 4'b1111;
        r_chickenpic[2690] <= 4'b1111;
        r_chickenpic[2691] <= 4'b1111;
        r_chickenpic[2692] <= 4'b1111;
        r_chickenpic[2693] <= 4'b1111;
        r_chickenpic[2694] <= 4'b1111;
        r_chickenpic[2695] <= 4'b1111;
        r_chickenpic[2696] <= 4'b1111;
        r_chickenpic[2697] <= 4'b1111;
        r_chickenpic[2698] <= 4'b1111;
        r_chickenpic[2699] <= 4'b1111;
        r_chickenpic[2700] <= 4'b1111;
        r_chickenpic[2701] <= 4'b1111;
        r_chickenpic[2702] <= 4'b1111;
        r_chickenpic[2703] <= 4'b1111;
        r_chickenpic[2704] <= 4'b1111;
        r_chickenpic[2705] <= 4'b1111;
        r_chickenpic[2706] <= 4'b1111;
        r_chickenpic[2707] <= 4'b1111;
        r_chickenpic[2708] <= 4'b1111;
        r_chickenpic[2709] <= 4'b1111;
        r_chickenpic[2710] <= 4'b1111;
        r_chickenpic[2711] <= 4'b1111;
        r_chickenpic[2712] <= 4'b1111;
        r_chickenpic[2713] <= 4'b1111;
        r_chickenpic[2714] <= 4'b1111;
        r_chickenpic[2715] <= 4'b1111;
        r_chickenpic[2716] <= 4'b1111;
        r_chickenpic[2717] <= 4'b1111;
        r_chickenpic[2718] <= 4'b1111;
        r_chickenpic[2719] <= 4'b1111;
        r_chickenpic[2720] <= 4'b1111;
        r_chickenpic[2721] <= 4'b1111;
        r_chickenpic[2722] <= 4'b1111;
        r_chickenpic[2723] <= 4'b1111;
        r_chickenpic[2724] <= 4'b0000;
        r_chickenpic[2725] <= 4'b0000;
        r_chickenpic[2726] <= 4'b0000;
        r_chickenpic[2727] <= 4'b1111;
        r_chickenpic[2728] <= 4'b1111;
        r_chickenpic[2729] <= 4'b1111;
        r_chickenpic[2730] <= 4'b1111;
        r_chickenpic[2731] <= 4'b1111;
        r_chickenpic[2732] <= 4'b1111;
        r_chickenpic[2733] <= 4'b1111;
        r_chickenpic[2734] <= 4'b1111;
        r_chickenpic[2735] <= 4'b1111;
        r_chickenpic[2736] <= 4'b1111;
        r_chickenpic[2737] <= 4'b1111;
        r_chickenpic[2738] <= 4'b1111;
        r_chickenpic[2739] <= 4'b1111;
        r_chickenpic[2740] <= 4'b1111;
        r_chickenpic[2741] <= 4'b1111;
        r_chickenpic[2742] <= 4'b1111;
        r_chickenpic[2743] <= 4'b1111;
        r_chickenpic[2744] <= 4'b1111;
        r_chickenpic[2745] <= 4'b1111;
        r_chickenpic[2746] <= 4'b1111;
        r_chickenpic[2747] <= 4'b1111;
        r_chickenpic[2748] <= 4'b1111;
        r_chickenpic[2749] <= 4'b1111;
        r_chickenpic[2750] <= 4'b1111;
        r_chickenpic[2751] <= 4'b1111;
        r_chickenpic[2752] <= 4'b1111;
        r_chickenpic[2753] <= 4'b1111;
        r_chickenpic[2754] <= 4'b1111;
        r_chickenpic[2755] <= 4'b1111;
        r_chickenpic[2756] <= 4'b1111;
        r_chickenpic[2757] <= 4'b1111;
        r_chickenpic[2758] <= 4'b1111;
        r_chickenpic[2759] <= 4'b1111;
        r_chickenpic[2760] <= 4'b1111;
        r_chickenpic[2761] <= 4'b1111;
        r_chickenpic[2762] <= 4'b1111;
        r_chickenpic[2763] <= 4'b1111;
        r_chickenpic[2764] <= 4'b1111;
        r_chickenpic[2765] <= 4'b1111;
        r_chickenpic[2766] <= 4'b1111;
        r_chickenpic[2767] <= 4'b1111;
        r_chickenpic[2768] <= 4'b1111;
        r_chickenpic[2769] <= 4'b1111;
        r_chickenpic[2770] <= 4'b1111;
        r_chickenpic[2771] <= 4'b1111;
        r_chickenpic[2772] <= 4'b1111;
        r_chickenpic[2773] <= 4'b1111;
        r_chickenpic[2774] <= 4'b1111;
        r_chickenpic[2775] <= 4'b1111;
        r_chickenpic[2776] <= 4'b1111;
        r_chickenpic[2777] <= 4'b1111;
        r_chickenpic[2778] <= 4'b0000;
        r_chickenpic[2779] <= 4'b0000;
        r_chickenpic[2780] <= 4'b1111;
        r_chickenpic[2781] <= 4'b1111;
        r_chickenpic[2782] <= 4'b1111;
        r_chickenpic[2783] <= 4'b1111;
        r_chickenpic[2784] <= 4'b1111;
        r_chickenpic[2785] <= 4'b1111;
        r_chickenpic[2786] <= 4'b1111;
        r_chickenpic[2787] <= 4'b1111;
        r_chickenpic[2788] <= 4'b1111;
        r_chickenpic[2789] <= 4'b1111;
        r_chickenpic[2790] <= 4'b1111;
        r_chickenpic[2791] <= 4'b1111;
        r_chickenpic[2792] <= 4'b1111;
        r_chickenpic[2793] <= 4'b1111;
        r_chickenpic[2794] <= 4'b1111;
        r_chickenpic[2795] <= 4'b1111;
        r_chickenpic[2796] <= 4'b1111;
        r_chickenpic[2797] <= 4'b1111;
        r_chickenpic[2798] <= 4'b1111;
        r_chickenpic[2799] <= 4'b1111;
        r_chickenpic[2800] <= 4'b1111;
        r_chickenpic[2801] <= 4'b1111;
        r_chickenpic[2802] <= 4'b1111;
        r_chickenpic[2803] <= 4'b1111;
        r_chickenpic[2804] <= 4'b1111;
        r_chickenpic[2805] <= 4'b1111;
        r_chickenpic[2806] <= 4'b1111;
        r_chickenpic[2807] <= 4'b1111;
        r_chickenpic[2808] <= 4'b1111;
        r_chickenpic[2809] <= 4'b1111;
        r_chickenpic[2810] <= 4'b1111;
        r_chickenpic[2811] <= 4'b1111;
        r_chickenpic[2812] <= 4'b1111;
        r_chickenpic[2813] <= 4'b1111;
        r_chickenpic[2814] <= 4'b1111;
        r_chickenpic[2815] <= 4'b1111;
        r_chickenpic[2816] <= 4'b1111;
        r_chickenpic[2817] <= 4'b1111;
        r_chickenpic[2818] <= 4'b1111;
        r_chickenpic[2819] <= 4'b1111;
        r_chickenpic[2820] <= 4'b1111;
        r_chickenpic[2821] <= 4'b1111;
        r_chickenpic[2822] <= 4'b1111;
        r_chickenpic[2823] <= 4'b1111;
        r_chickenpic[2824] <= 4'b1111;
        r_chickenpic[2825] <= 4'b1111;
        r_chickenpic[2826] <= 4'b1111;
        r_chickenpic[2827] <= 4'b1111;
        r_chickenpic[2828] <= 4'b1111;
        r_chickenpic[2829] <= 4'b1111;
        r_chickenpic[2830] <= 4'b1111;
        r_chickenpic[2831] <= 4'b1111;
        r_chickenpic[2832] <= 4'b1111;
        r_chickenpic[2833] <= 4'b1111;
        r_chickenpic[2834] <= 4'b1111;
        r_chickenpic[2835] <= 4'b1111;
        r_chickenpic[2836] <= 4'b1111;
        r_chickenpic[2837] <= 4'b1111;
        r_chickenpic[2838] <= 4'b1111;
        r_chickenpic[2839] <= 4'b1111;
        r_chickenpic[2840] <= 4'b1111;
        r_chickenpic[2841] <= 4'b1111;
        r_chickenpic[2842] <= 4'b1111;
        r_chickenpic[2843] <= 4'b1111;
        r_chickenpic[2844] <= 4'b1111;
        r_chickenpic[2845] <= 4'b1111;
        r_chickenpic[2846] <= 4'b1111;
        r_chickenpic[2847] <= 4'b1111;
        r_chickenpic[2848] <= 4'b1111;
        r_chickenpic[2849] <= 4'b1111;
        r_chickenpic[2850] <= 4'b1111;
        r_chickenpic[2851] <= 4'b1111;
        r_chickenpic[2852] <= 4'b1111;
        r_chickenpic[2853] <= 4'b1111;
        r_chickenpic[2854] <= 4'b1111;
        r_chickenpic[2855] <= 4'b1111;
        r_chickenpic[2856] <= 4'b1111;
        r_chickenpic[2857] <= 4'b1111;
        r_chickenpic[2858] <= 4'b1111;
        r_chickenpic[2859] <= 4'b1111;
        r_chickenpic[2860] <= 4'b1111;
        r_chickenpic[2861] <= 4'b1111;
        r_chickenpic[2862] <= 4'b1111;
        r_chickenpic[2863] <= 4'b1111;
        r_chickenpic[2864] <= 4'b1111;
        r_chickenpic[2865] <= 4'b1111;
        r_chickenpic[2866] <= 4'b1111;
        r_chickenpic[2867] <= 4'b1111;
        r_chickenpic[2868] <= 4'b1111;
        r_chickenpic[2869] <= 4'b1111;
        r_chickenpic[2870] <= 4'b1111;
        r_chickenpic[2871] <= 4'b1111;
        r_chickenpic[2872] <= 4'b1111;
        r_chickenpic[2873] <= 4'b1111;
        r_chickenpic[2874] <= 4'b1111;
        r_chickenpic[2875] <= 4'b1111;
        r_chickenpic[2876] <= 4'b1111;
        r_chickenpic[2877] <= 4'b1111;
        r_chickenpic[2878] <= 4'b1111;
        r_chickenpic[2879] <= 4'b1111;
        r_chickenpic[2880] <= 4'b1111;
        r_chickenpic[2881] <= 4'b1111;
        r_chickenpic[2882] <= 4'b1111;
        r_chickenpic[2883] <= 4'b1111;
        r_chickenpic[2884] <= 4'b1111;
        r_chickenpic[2885] <= 4'b1111;
        r_chickenpic[2886] <= 4'b1111;
        r_chickenpic[2887] <= 4'b1111;
        r_chickenpic[2888] <= 4'b1111;
        r_chickenpic[2889] <= 4'b1111;
        r_chickenpic[2890] <= 4'b1111;
        r_chickenpic[2891] <= 4'b1111;
        r_chickenpic[2892] <= 4'b1111;
        r_chickenpic[2893] <= 4'b1111;
        r_chickenpic[2894] <= 4'b1111;
        r_chickenpic[2895] <= 4'b1111;
        r_chickenpic[2896] <= 4'b1111;
        r_chickenpic[2897] <= 4'b1111;
        r_chickenpic[2898] <= 4'b1111;
        r_chickenpic[2899] <= 4'b1111;
        r_chickenpic[2900] <= 4'b1111;
        r_chickenpic[2901] <= 4'b1111;
        r_chickenpic[2902] <= 4'b1111;
        r_chickenpic[2903] <= 4'b1111;
        r_chickenpic[2904] <= 4'b1111;
        r_chickenpic[2905] <= 4'b1111;
        r_chickenpic[2906] <= 4'b1111;
        r_chickenpic[2907] <= 4'b1111;
        r_chickenpic[2908] <= 4'b1111;
        r_chickenpic[2909] <= 4'b1111;
        r_chickenpic[2910] <= 4'b1111;
        r_chickenpic[2911] <= 4'b1111;
        r_chickenpic[2912] <= 4'b1111;
        r_chickenpic[2913] <= 4'b1111;
        r_chickenpic[2914] <= 4'b1111;
        r_chickenpic[2915] <= 4'b1111;
        r_chickenpic[2916] <= 4'b1111;
        r_chickenpic[2917] <= 4'b1111;
        r_chickenpic[2918] <= 4'b1111;
        r_chickenpic[2919] <= 4'b1111;
        r_chickenpic[2920] <= 4'b1111;
        r_chickenpic[2921] <= 4'b1111;
        r_chickenpic[2922] <= 4'b1111;
        r_chickenpic[2923] <= 4'b1111;
        r_chickenpic[2924] <= 4'b1111;
        r_chickenpic[2925] <= 4'b1111;
        r_chickenpic[2926] <= 4'b1111;
        r_chickenpic[2927] <= 4'b1111;
        r_chickenpic[2928] <= 4'b1111;
        r_chickenpic[2929] <= 4'b1111;
        r_chickenpic[2930] <= 4'b1111;
        r_chickenpic[2931] <= 4'b1111;
        r_chickenpic[2932] <= 4'b1111;
        r_chickenpic[2933] <= 4'b1111;
        r_chickenpic[2934] <= 4'b1111;
        r_chickenpic[2935] <= 4'b1111;
        r_chickenpic[2936] <= 4'b1111;
        r_chickenpic[2937] <= 4'b1111;
        r_chickenpic[2938] <= 4'b1111;
        r_chickenpic[2939] <= 4'b1111;
        r_chickenpic[2940] <= 4'b1111;
        r_chickenpic[2941] <= 4'b1111;
        r_chickenpic[2942] <= 4'b1111;
        r_chickenpic[2943] <= 4'b1111;
        r_chickenpic[2944] <= 4'b1111;
        r_chickenpic[2945] <= 4'b1111;
        r_chickenpic[2946] <= 4'b1111;
        r_chickenpic[2947] <= 4'b1111;
        r_chickenpic[2948] <= 4'b1111;
        r_chickenpic[2949] <= 4'b1111;
        r_chickenpic[2950] <= 4'b1111;
        r_chickenpic[2951] <= 4'b1111;
        r_chickenpic[2952] <= 4'b1111;
        r_chickenpic[2953] <= 4'b1111;
        r_chickenpic[2954] <= 4'b1111;
        r_chickenpic[2955] <= 4'b1111;
        r_chickenpic[2956] <= 4'b1111;
        r_chickenpic[2957] <= 4'b1111;
        r_chickenpic[2958] <= 4'b1111;
        r_chickenpic[2959] <= 4'b1111;
        r_chickenpic[2960] <= 4'b1111;
        r_chickenpic[2961] <= 4'b1111;
        r_chickenpic[2962] <= 4'b1111;
        r_chickenpic[2963] <= 4'b1111;
        r_chickenpic[2964] <= 4'b1111;
        r_chickenpic[2965] <= 4'b1111;
        r_chickenpic[2966] <= 4'b1111;
        r_chickenpic[2967] <= 4'b1111;
        r_chickenpic[2968] <= 4'b1111;
        r_chickenpic[2969] <= 4'b1111;
        r_chickenpic[2970] <= 4'b1111;
        r_chickenpic[2971] <= 4'b1111;
        r_chickenpic[2972] <= 4'b1111;
        r_chickenpic[2973] <= 4'b1111;
        r_chickenpic[2974] <= 4'b1111;
        r_chickenpic[2975] <= 4'b1111;
        r_chickenpic[2976] <= 4'b1111;
        r_chickenpic[2977] <= 4'b1111;
        r_chickenpic[2978] <= 4'b1111;
        r_chickenpic[2979] <= 4'b1111;
        r_chickenpic[2980] <= 4'b1111;
        r_chickenpic[2981] <= 4'b1111;
        r_chickenpic[2982] <= 4'b1111;
        r_chickenpic[2983] <= 4'b1111;
        r_chickenpic[2984] <= 4'b1111;
        r_chickenpic[2985] <= 4'b1111;
        r_chickenpic[2986] <= 4'b1111;
        r_chickenpic[2987] <= 4'b1111;
        r_chickenpic[2988] <= 4'b1111;
        r_chickenpic[2989] <= 4'b1111;
        r_chickenpic[2990] <= 4'b1111;
        r_chickenpic[2991] <= 4'b1111;
        r_chickenpic[2992] <= 4'b1111;
        r_chickenpic[2993] <= 4'b1111;
        r_chickenpic[2994] <= 4'b1111;
        r_chickenpic[2995] <= 4'b1111;
        r_chickenpic[2996] <= 4'b1111;
        r_chickenpic[2997] <= 4'b1111;
        r_chickenpic[2998] <= 4'b1111;
        r_chickenpic[2999] <= 4'b1111;
        r_chickenpic[3000] <= 4'b1111;
        r_chickenpic[3001] <= 4'b1111;
        r_chickenpic[3002] <= 4'b1111;
        r_chickenpic[3003] <= 4'b1111;
        r_chickenpic[3004] <= 4'b1111;
        r_chickenpic[3005] <= 4'b1111;
        r_chickenpic[3006] <= 4'b1111;
        r_chickenpic[3007] <= 4'b1111;
        r_chickenpic[3008] <= 4'b1111;
        r_chickenpic[3009] <= 4'b1111;
        r_chickenpic[3010] <= 4'b1111;
        r_chickenpic[3011] <= 4'b1111;
        r_chickenpic[3012] <= 4'b1111;
        r_chickenpic[3013] <= 4'b1111;
        r_chickenpic[3014] <= 4'b1111;
        r_chickenpic[3015] <= 4'b1111;
        r_chickenpic[3016] <= 4'b1111;
        r_chickenpic[3017] <= 4'b1111;
        r_chickenpic[3018] <= 4'b1111;
        r_chickenpic[3019] <= 4'b1111;
        r_chickenpic[3020] <= 4'b1111;
        r_chickenpic[3021] <= 4'b1111;
        r_chickenpic[3022] <= 4'b1111;
        r_chickenpic[3023] <= 4'b1111;
        r_chickenpic[3024] <= 4'b1111;

        r_rabbitpic[0] <= 4'b1111;
        r_rabbitpic[1] <= 4'b1111;
        r_rabbitpic[2] <= 4'b1111;
        r_rabbitpic[3] <= 4'b1111;
        r_rabbitpic[4] <= 4'b1111;
        r_rabbitpic[5] <= 4'b1111;
        r_rabbitpic[6] <= 4'b1111;
        r_rabbitpic[7] <= 4'b1111;
        r_rabbitpic[8] <= 4'b1111;
        r_rabbitpic[9] <= 4'b1111;
        r_rabbitpic[10] <= 4'b1111;
        r_rabbitpic[11] <= 4'b1111;
        r_rabbitpic[12] <= 4'b1111;
        r_rabbitpic[13] <= 4'b1111;
        r_rabbitpic[14] <= 4'b1111;
        r_rabbitpic[15] <= 4'b1111;
        r_rabbitpic[16] <= 4'b1111;
        r_rabbitpic[17] <= 4'b1111;
        r_rabbitpic[18] <= 4'b1111;
        r_rabbitpic[19] <= 4'b1111;
        r_rabbitpic[20] <= 4'b1111;
        r_rabbitpic[21] <= 4'b1111;
        r_rabbitpic[22] <= 4'b1111;
        r_rabbitpic[23] <= 4'b1111;
        r_rabbitpic[24] <= 4'b1111;
        r_rabbitpic[25] <= 4'b1111;
        r_rabbitpic[26] <= 4'b1111;
        r_rabbitpic[27] <= 4'b1111;
        r_rabbitpic[28] <= 4'b1111;
        r_rabbitpic[29] <= 4'b1111;
        r_rabbitpic[30] <= 4'b1111;
        r_rabbitpic[31] <= 4'b1111;
        r_rabbitpic[32] <= 4'b1111;
        r_rabbitpic[33] <= 4'b1111;
        r_rabbitpic[34] <= 4'b1111;
        r_rabbitpic[35] <= 4'b1111;
        r_rabbitpic[36] <= 4'b1111;
        r_rabbitpic[37] <= 4'b1111;
        r_rabbitpic[38] <= 4'b1111;
        r_rabbitpic[39] <= 4'b1111;
        r_rabbitpic[40] <= 4'b1111;
        r_rabbitpic[41] <= 4'b1111;
        r_rabbitpic[42] <= 4'b1111;
        r_rabbitpic[43] <= 4'b1111;
        r_rabbitpic[44] <= 4'b1111;
        r_rabbitpic[45] <= 4'b1111;
        r_rabbitpic[46] <= 4'b1111;
        r_rabbitpic[47] <= 4'b1111;
        r_rabbitpic[48] <= 4'b1111;
        r_rabbitpic[49] <= 4'b1111;
        r_rabbitpic[50] <= 4'b1111;
        r_rabbitpic[51] <= 4'b1111;
        r_rabbitpic[52] <= 4'b1111;
        r_rabbitpic[53] <= 4'b1111;
        r_rabbitpic[54] <= 4'b1111;
        r_rabbitpic[55] <= 4'b1111;
        r_rabbitpic[56] <= 4'b1111;
        r_rabbitpic[57] <= 4'b1111;
        r_rabbitpic[58] <= 4'b1111;
        r_rabbitpic[59] <= 4'b1111;
        r_rabbitpic[60] <= 4'b1111;
        r_rabbitpic[61] <= 4'b1111;
        r_rabbitpic[62] <= 4'b1111;
        r_rabbitpic[63] <= 4'b1111;
        r_rabbitpic[64] <= 4'b1111;
        r_rabbitpic[65] <= 4'b1111;
        r_rabbitpic[66] <= 4'b1111;
        r_rabbitpic[67] <= 4'b1111;
        r_rabbitpic[68] <= 4'b1111;
        r_rabbitpic[69] <= 4'b1111;
        r_rabbitpic[70] <= 4'b1111;
        r_rabbitpic[71] <= 4'b1111;
        r_rabbitpic[72] <= 4'b1111;
        r_rabbitpic[73] <= 4'b1111;
        r_rabbitpic[74] <= 4'b1111;
        r_rabbitpic[75] <= 4'b1111;
        r_rabbitpic[76] <= 4'b1111;
        r_rabbitpic[77] <= 4'b1111;
        r_rabbitpic[78] <= 4'b1111;
        r_rabbitpic[79] <= 4'b1111;
        r_rabbitpic[80] <= 4'b1111;
        r_rabbitpic[81] <= 4'b1111;
        r_rabbitpic[82] <= 4'b1111;
        r_rabbitpic[83] <= 4'b1111;
        r_rabbitpic[84] <= 4'b1111;
        r_rabbitpic[85] <= 4'b1111;
        r_rabbitpic[86] <= 4'b1111;
        r_rabbitpic[87] <= 4'b1111;
        r_rabbitpic[88] <= 4'b1111;
        r_rabbitpic[89] <= 4'b1111;
        r_rabbitpic[90] <= 4'b1111;
        r_rabbitpic[91] <= 4'b1111;
        r_rabbitpic[92] <= 4'b1111;
        r_rabbitpic[93] <= 4'b1111;
        r_rabbitpic[94] <= 4'b1111;
        r_rabbitpic[95] <= 4'b1111;
        r_rabbitpic[96] <= 4'b1111;
        r_rabbitpic[97] <= 4'b1111;
        r_rabbitpic[98] <= 4'b1111;
        r_rabbitpic[99] <= 4'b1111;
        r_rabbitpic[100] <= 4'b1111;
        r_rabbitpic[101] <= 4'b1111;
        r_rabbitpic[102] <= 4'b1111;
        r_rabbitpic[103] <= 4'b1111;
        r_rabbitpic[104] <= 4'b1111;
        r_rabbitpic[105] <= 4'b1111;
        r_rabbitpic[106] <= 4'b1111;
        r_rabbitpic[107] <= 4'b1111;
        r_rabbitpic[108] <= 4'b1111;
        r_rabbitpic[109] <= 4'b1111;
        r_rabbitpic[110] <= 4'b1111;
        r_rabbitpic[111] <= 4'b1111;
        r_rabbitpic[112] <= 4'b1111;
        r_rabbitpic[113] <= 4'b1111;
        r_rabbitpic[114] <= 4'b1111;
        r_rabbitpic[115] <= 4'b1111;
        r_rabbitpic[116] <= 4'b1111;
        r_rabbitpic[117] <= 4'b1111;
        r_rabbitpic[118] <= 4'b1111;
        r_rabbitpic[119] <= 4'b1111;
        r_rabbitpic[120] <= 4'b1111;
        r_rabbitpic[121] <= 4'b1111;
        r_rabbitpic[122] <= 4'b1111;
        r_rabbitpic[123] <= 4'b1111;
        r_rabbitpic[124] <= 4'b1111;
        r_rabbitpic[125] <= 4'b1111;
        r_rabbitpic[126] <= 4'b1111;
        r_rabbitpic[127] <= 4'b1111;
        r_rabbitpic[128] <= 4'b1111;
        r_rabbitpic[129] <= 4'b1111;
        r_rabbitpic[130] <= 4'b1111;
        r_rabbitpic[131] <= 4'b1111;
        r_rabbitpic[132] <= 4'b1111;
        r_rabbitpic[133] <= 4'b1111;
        r_rabbitpic[134] <= 4'b1111;
        r_rabbitpic[135] <= 4'b1111;
        r_rabbitpic[136] <= 4'b1111;
        r_rabbitpic[137] <= 4'b1111;
        r_rabbitpic[138] <= 4'b1111;
        r_rabbitpic[139] <= 4'b1111;
        r_rabbitpic[140] <= 4'b1111;
        r_rabbitpic[141] <= 4'b1111;
        r_rabbitpic[142] <= 4'b1111;
        r_rabbitpic[143] <= 4'b1111;
        r_rabbitpic[144] <= 4'b1111;
        r_rabbitpic[145] <= 4'b1111;
        r_rabbitpic[146] <= 4'b1111;
        r_rabbitpic[147] <= 4'b1111;
        r_rabbitpic[148] <= 4'b1111;
        r_rabbitpic[149] <= 4'b1111;
        r_rabbitpic[150] <= 4'b1111;
        r_rabbitpic[151] <= 4'b1111;
        r_rabbitpic[152] <= 4'b1111;
        r_rabbitpic[153] <= 4'b1111;
        r_rabbitpic[154] <= 4'b1111;
        r_rabbitpic[155] <= 4'b1111;
        r_rabbitpic[156] <= 4'b1111;
        r_rabbitpic[157] <= 4'b1111;
        r_rabbitpic[158] <= 4'b1111;
        r_rabbitpic[159] <= 4'b1111;
        r_rabbitpic[160] <= 4'b1111;
        r_rabbitpic[161] <= 4'b1111;
        r_rabbitpic[162] <= 4'b1111;
        r_rabbitpic[163] <= 4'b1111;
        r_rabbitpic[164] <= 4'b1111;
        r_rabbitpic[165] <= 4'b1111;
        r_rabbitpic[166] <= 4'b1111;
        r_rabbitpic[167] <= 4'b1111;
        r_rabbitpic[168] <= 4'b1111;
        r_rabbitpic[169] <= 4'b1111;
        r_rabbitpic[170] <= 4'b1111;
        r_rabbitpic[171] <= 4'b1111;
        r_rabbitpic[172] <= 4'b1111;
        r_rabbitpic[173] <= 4'b1111;
        r_rabbitpic[174] <= 4'b1111;
        r_rabbitpic[175] <= 4'b1111;
        r_rabbitpic[176] <= 4'b1111;
        r_rabbitpic[177] <= 4'b1111;
        r_rabbitpic[178] <= 4'b1111;
        r_rabbitpic[179] <= 4'b1111;
        r_rabbitpic[180] <= 4'b1111;
        r_rabbitpic[181] <= 4'b1111;
        r_rabbitpic[182] <= 4'b1111;
        r_rabbitpic[183] <= 4'b1111;
        r_rabbitpic[184] <= 4'b1111;
        r_rabbitpic[185] <= 4'b1111;
        r_rabbitpic[186] <= 4'b1111;
        r_rabbitpic[187] <= 4'b1111;
        r_rabbitpic[188] <= 4'b1111;
        r_rabbitpic[189] <= 4'b1111;
        r_rabbitpic[190] <= 4'b1111;
        r_rabbitpic[191] <= 4'b1111;
        r_rabbitpic[192] <= 4'b1111;
        r_rabbitpic[193] <= 4'b1111;
        r_rabbitpic[194] <= 4'b1111;
        r_rabbitpic[195] <= 4'b1111;
        r_rabbitpic[196] <= 4'b1111;
        r_rabbitpic[197] <= 4'b1111;
        r_rabbitpic[198] <= 4'b1111;
        r_rabbitpic[199] <= 4'b1111;
        r_rabbitpic[200] <= 4'b1111;
        r_rabbitpic[201] <= 4'b1111;
        r_rabbitpic[202] <= 4'b1111;
        r_rabbitpic[203] <= 4'b1111;
        r_rabbitpic[204] <= 4'b1111;
        r_rabbitpic[205] <= 4'b1111;
        r_rabbitpic[206] <= 4'b1111;
        r_rabbitpic[207] <= 4'b1111;
        r_rabbitpic[208] <= 4'b1111;
        r_rabbitpic[209] <= 4'b1111;
        r_rabbitpic[210] <= 4'b1111;
        r_rabbitpic[211] <= 4'b1111;
        r_rabbitpic[212] <= 4'b1111;
        r_rabbitpic[213] <= 4'b1111;
        r_rabbitpic[214] <= 4'b1111;
        r_rabbitpic[215] <= 4'b1111;
        r_rabbitpic[216] <= 4'b1111;
        r_rabbitpic[217] <= 4'b1111;
        r_rabbitpic[218] <= 4'b1111;
        r_rabbitpic[219] <= 4'b1111;
        r_rabbitpic[220] <= 4'b1111;
        r_rabbitpic[221] <= 4'b1111;
        r_rabbitpic[222] <= 4'b1111;
        r_rabbitpic[223] <= 4'b1111;
        r_rabbitpic[224] <= 4'b1111;
        r_rabbitpic[225] <= 4'b1111;
        r_rabbitpic[226] <= 4'b1111;
        r_rabbitpic[227] <= 4'b1111;
        r_rabbitpic[228] <= 4'b1111;
        r_rabbitpic[229] <= 4'b1111;
        r_rabbitpic[230] <= 4'b1111;
        r_rabbitpic[231] <= 4'b1111;
        r_rabbitpic[232] <= 4'b1111;
        r_rabbitpic[233] <= 4'b1111;
        r_rabbitpic[234] <= 4'b1111;
        r_rabbitpic[235] <= 4'b1111;
        r_rabbitpic[236] <= 4'b0000;
        r_rabbitpic[237] <= 4'b0000;
        r_rabbitpic[238] <= 4'b1111;
        r_rabbitpic[239] <= 4'b1111;
        r_rabbitpic[240] <= 4'b1111;
        r_rabbitpic[241] <= 4'b1111;
        r_rabbitpic[242] <= 4'b1111;
        r_rabbitpic[243] <= 4'b1111;
        r_rabbitpic[244] <= 4'b1111;
        r_rabbitpic[245] <= 4'b1111;
        r_rabbitpic[246] <= 4'b0000;
        r_rabbitpic[247] <= 4'b0000;
        r_rabbitpic[248] <= 4'b1111;
        r_rabbitpic[249] <= 4'b1111;
        r_rabbitpic[250] <= 4'b1111;
        r_rabbitpic[251] <= 4'b1111;
        r_rabbitpic[252] <= 4'b1111;
        r_rabbitpic[253] <= 4'b1111;
        r_rabbitpic[254] <= 4'b1111;
        r_rabbitpic[255] <= 4'b1111;
        r_rabbitpic[256] <= 4'b1111;
        r_rabbitpic[257] <= 4'b1111;
        r_rabbitpic[258] <= 4'b1111;
        r_rabbitpic[259] <= 4'b1111;
        r_rabbitpic[260] <= 4'b1111;
        r_rabbitpic[261] <= 4'b1111;
        r_rabbitpic[262] <= 4'b1111;
        r_rabbitpic[263] <= 4'b1111;
        r_rabbitpic[264] <= 4'b1111;
        r_rabbitpic[265] <= 4'b1111;
        r_rabbitpic[266] <= 4'b1111;
        r_rabbitpic[267] <= 4'b1111;
        r_rabbitpic[268] <= 4'b1111;
        r_rabbitpic[269] <= 4'b1111;
        r_rabbitpic[270] <= 4'b1111;
        r_rabbitpic[271] <= 4'b1111;
        r_rabbitpic[272] <= 4'b1111;
        r_rabbitpic[273] <= 4'b1111;
        r_rabbitpic[274] <= 4'b1111;
        r_rabbitpic[275] <= 4'b1111;
        r_rabbitpic[276] <= 4'b1111;
        r_rabbitpic[277] <= 4'b1111;
        r_rabbitpic[278] <= 4'b1111;
        r_rabbitpic[279] <= 4'b1111;
        r_rabbitpic[280] <= 4'b1111;
        r_rabbitpic[281] <= 4'b1111;
        r_rabbitpic[282] <= 4'b1111;
        r_rabbitpic[283] <= 4'b1111;
        r_rabbitpic[284] <= 4'b1111;
        r_rabbitpic[285] <= 4'b1111;
        r_rabbitpic[286] <= 4'b1111;
        r_rabbitpic[287] <= 4'b1111;
        r_rabbitpic[288] <= 4'b1111;
        r_rabbitpic[289] <= 4'b1111;
        r_rabbitpic[290] <= 4'b0000;
        r_rabbitpic[291] <= 4'b1111;
        r_rabbitpic[292] <= 4'b0000;
        r_rabbitpic[293] <= 4'b0000;
        r_rabbitpic[294] <= 4'b1111;
        r_rabbitpic[295] <= 4'b1111;
        r_rabbitpic[296] <= 4'b1111;
        r_rabbitpic[297] <= 4'b1111;
        r_rabbitpic[298] <= 4'b1111;
        r_rabbitpic[299] <= 4'b1111;
        r_rabbitpic[300] <= 4'b0000;
        r_rabbitpic[301] <= 4'b0000;
        r_rabbitpic[302] <= 4'b1111;
        r_rabbitpic[303] <= 4'b1111;
        r_rabbitpic[304] <= 4'b1111;
        r_rabbitpic[305] <= 4'b1111;
        r_rabbitpic[306] <= 4'b1111;
        r_rabbitpic[307] <= 4'b1111;
        r_rabbitpic[308] <= 4'b1111;
        r_rabbitpic[309] <= 4'b1111;
        r_rabbitpic[310] <= 4'b1111;
        r_rabbitpic[311] <= 4'b1111;
        r_rabbitpic[312] <= 4'b1111;
        r_rabbitpic[313] <= 4'b1111;
        r_rabbitpic[314] <= 4'b1111;
        r_rabbitpic[315] <= 4'b1111;
        r_rabbitpic[316] <= 4'b1111;
        r_rabbitpic[317] <= 4'b1111;
        r_rabbitpic[318] <= 4'b1111;
        r_rabbitpic[319] <= 4'b1111;
        r_rabbitpic[320] <= 4'b1111;
        r_rabbitpic[321] <= 4'b1111;
        r_rabbitpic[322] <= 4'b1111;
        r_rabbitpic[323] <= 4'b1111;
        r_rabbitpic[324] <= 4'b1111;
        r_rabbitpic[325] <= 4'b1111;
        r_rabbitpic[326] <= 4'b1111;
        r_rabbitpic[327] <= 4'b1111;
        r_rabbitpic[328] <= 4'b1111;
        r_rabbitpic[329] <= 4'b1111;
        r_rabbitpic[330] <= 4'b1111;
        r_rabbitpic[331] <= 4'b1111;
        r_rabbitpic[332] <= 4'b1111;
        r_rabbitpic[333] <= 4'b1111;
        r_rabbitpic[334] <= 4'b1111;
        r_rabbitpic[335] <= 4'b1111;
        r_rabbitpic[336] <= 4'b1111;
        r_rabbitpic[337] <= 4'b1111;
        r_rabbitpic[338] <= 4'b1111;
        r_rabbitpic[339] <= 4'b1111;
        r_rabbitpic[340] <= 4'b1111;
        r_rabbitpic[341] <= 4'b1111;
        r_rabbitpic[342] <= 4'b1111;
        r_rabbitpic[343] <= 4'b1111;
        r_rabbitpic[344] <= 4'b1111;
        r_rabbitpic[345] <= 4'b1111;
        r_rabbitpic[346] <= 4'b1111;
        r_rabbitpic[347] <= 4'b1111;
        r_rabbitpic[348] <= 4'b0000;
        r_rabbitpic[349] <= 4'b1111;
        r_rabbitpic[350] <= 4'b1111;
        r_rabbitpic[351] <= 4'b1111;
        r_rabbitpic[352] <= 4'b1111;
        r_rabbitpic[353] <= 4'b1111;
        r_rabbitpic[354] <= 4'b1111;
        r_rabbitpic[355] <= 4'b0000;
        r_rabbitpic[356] <= 4'b1111;
        r_rabbitpic[357] <= 4'b1111;
        r_rabbitpic[358] <= 4'b1111;
        r_rabbitpic[359] <= 4'b1111;
        r_rabbitpic[360] <= 4'b1111;
        r_rabbitpic[361] <= 4'b1111;
        r_rabbitpic[362] <= 4'b1111;
        r_rabbitpic[363] <= 4'b1111;
        r_rabbitpic[364] <= 4'b1111;
        r_rabbitpic[365] <= 4'b1111;
        r_rabbitpic[366] <= 4'b1111;
        r_rabbitpic[367] <= 4'b1111;
        r_rabbitpic[368] <= 4'b1111;
        r_rabbitpic[369] <= 4'b1111;
        r_rabbitpic[370] <= 4'b1111;
        r_rabbitpic[371] <= 4'b1111;
        r_rabbitpic[372] <= 4'b1111;
        r_rabbitpic[373] <= 4'b1111;
        r_rabbitpic[374] <= 4'b1111;
        r_rabbitpic[375] <= 4'b1111;
        r_rabbitpic[376] <= 4'b1111;
        r_rabbitpic[377] <= 4'b1111;
        r_rabbitpic[378] <= 4'b1111;
        r_rabbitpic[379] <= 4'b1111;
        r_rabbitpic[380] <= 4'b1111;
        r_rabbitpic[381] <= 4'b1111;
        r_rabbitpic[382] <= 4'b1111;
        r_rabbitpic[383] <= 4'b1111;
        r_rabbitpic[384] <= 4'b1111;
        r_rabbitpic[385] <= 4'b1111;
        r_rabbitpic[386] <= 4'b1111;
        r_rabbitpic[387] <= 4'b1111;
        r_rabbitpic[388] <= 4'b1111;
        r_rabbitpic[389] <= 4'b1111;
        r_rabbitpic[390] <= 4'b1111;
        r_rabbitpic[391] <= 4'b1111;
        r_rabbitpic[392] <= 4'b1111;
        r_rabbitpic[393] <= 4'b1111;
        r_rabbitpic[394] <= 4'b1111;
        r_rabbitpic[395] <= 4'b1111;
        r_rabbitpic[396] <= 4'b1111;
        r_rabbitpic[397] <= 4'b1111;
        r_rabbitpic[398] <= 4'b1111;
        r_rabbitpic[399] <= 4'b1111;
        r_rabbitpic[400] <= 4'b1111;
        r_rabbitpic[401] <= 4'b0000;
        r_rabbitpic[402] <= 4'b1111;
        r_rabbitpic[403] <= 4'b0000;
        r_rabbitpic[404] <= 4'b0000;
        r_rabbitpic[405] <= 4'b1111;
        r_rabbitpic[406] <= 4'b1111;
        r_rabbitpic[407] <= 4'b1111;
        r_rabbitpic[408] <= 4'b1111;
        r_rabbitpic[409] <= 4'b0000;
        r_rabbitpic[410] <= 4'b0000;
        r_rabbitpic[411] <= 4'b1111;
        r_rabbitpic[412] <= 4'b0000;
        r_rabbitpic[413] <= 4'b1111;
        r_rabbitpic[414] <= 4'b1111;
        r_rabbitpic[415] <= 4'b1111;
        r_rabbitpic[416] <= 4'b1111;
        r_rabbitpic[417] <= 4'b1111;
        r_rabbitpic[418] <= 4'b1111;
        r_rabbitpic[419] <= 4'b1111;
        r_rabbitpic[420] <= 4'b1111;
        r_rabbitpic[421] <= 4'b1111;
        r_rabbitpic[422] <= 4'b1111;
        r_rabbitpic[423] <= 4'b1111;
        r_rabbitpic[424] <= 4'b1111;
        r_rabbitpic[425] <= 4'b1111;
        r_rabbitpic[426] <= 4'b1111;
        r_rabbitpic[427] <= 4'b1111;
        r_rabbitpic[428] <= 4'b1111;
        r_rabbitpic[429] <= 4'b1111;
        r_rabbitpic[430] <= 4'b1111;
        r_rabbitpic[431] <= 4'b1111;
        r_rabbitpic[432] <= 4'b1111;
        r_rabbitpic[433] <= 4'b1111;
        r_rabbitpic[434] <= 4'b1111;
        r_rabbitpic[435] <= 4'b1111;
        r_rabbitpic[436] <= 4'b1111;
        r_rabbitpic[437] <= 4'b1111;
        r_rabbitpic[438] <= 4'b1111;
        r_rabbitpic[439] <= 4'b1111;
        r_rabbitpic[440] <= 4'b1111;
        r_rabbitpic[441] <= 4'b1111;
        r_rabbitpic[442] <= 4'b1111;
        r_rabbitpic[443] <= 4'b1111;
        r_rabbitpic[444] <= 4'b1111;
        r_rabbitpic[445] <= 4'b1111;
        r_rabbitpic[446] <= 4'b1111;
        r_rabbitpic[447] <= 4'b1111;
        r_rabbitpic[448] <= 4'b1111;
        r_rabbitpic[449] <= 4'b1111;
        r_rabbitpic[450] <= 4'b1111;
        r_rabbitpic[451] <= 4'b1111;
        r_rabbitpic[452] <= 4'b1111;
        r_rabbitpic[453] <= 4'b1111;
        r_rabbitpic[454] <= 4'b1111;
        r_rabbitpic[455] <= 4'b1111;
        r_rabbitpic[456] <= 4'b0000;
        r_rabbitpic[457] <= 4'b1111;
        r_rabbitpic[458] <= 4'b1111;
        r_rabbitpic[459] <= 4'b0000;
        r_rabbitpic[460] <= 4'b0000;
        r_rabbitpic[461] <= 4'b1111;
        r_rabbitpic[462] <= 4'b1111;
        r_rabbitpic[463] <= 4'b0000;
        r_rabbitpic[464] <= 4'b0000;
        r_rabbitpic[465] <= 4'b1111;
        r_rabbitpic[466] <= 4'b1111;
        r_rabbitpic[467] <= 4'b0000;
        r_rabbitpic[468] <= 4'b1111;
        r_rabbitpic[469] <= 4'b1111;
        r_rabbitpic[470] <= 4'b1111;
        r_rabbitpic[471] <= 4'b1111;
        r_rabbitpic[472] <= 4'b1111;
        r_rabbitpic[473] <= 4'b1111;
        r_rabbitpic[474] <= 4'b1111;
        r_rabbitpic[475] <= 4'b1111;
        r_rabbitpic[476] <= 4'b1111;
        r_rabbitpic[477] <= 4'b1111;
        r_rabbitpic[478] <= 4'b1111;
        r_rabbitpic[479] <= 4'b1111;
        r_rabbitpic[480] <= 4'b1111;
        r_rabbitpic[481] <= 4'b1111;
        r_rabbitpic[482] <= 4'b1111;
        r_rabbitpic[483] <= 4'b1111;
        r_rabbitpic[484] <= 4'b1111;
        r_rabbitpic[485] <= 4'b1111;
        r_rabbitpic[486] <= 4'b1111;
        r_rabbitpic[487] <= 4'b1111;
        r_rabbitpic[488] <= 4'b1111;
        r_rabbitpic[489] <= 4'b1111;
        r_rabbitpic[490] <= 4'b1111;
        r_rabbitpic[491] <= 4'b1111;
        r_rabbitpic[492] <= 4'b1111;
        r_rabbitpic[493] <= 4'b1111;
        r_rabbitpic[494] <= 4'b1111;
        r_rabbitpic[495] <= 4'b1111;
        r_rabbitpic[496] <= 4'b1111;
        r_rabbitpic[497] <= 4'b1111;
        r_rabbitpic[498] <= 4'b1111;
        r_rabbitpic[499] <= 4'b1111;
        r_rabbitpic[500] <= 4'b1111;
        r_rabbitpic[501] <= 4'b1111;
        r_rabbitpic[502] <= 4'b1111;
        r_rabbitpic[503] <= 4'b1111;
        r_rabbitpic[504] <= 4'b1111;
        r_rabbitpic[505] <= 4'b1111;
        r_rabbitpic[506] <= 4'b1111;
        r_rabbitpic[507] <= 4'b1111;
        r_rabbitpic[508] <= 4'b1111;
        r_rabbitpic[509] <= 4'b1111;
        r_rabbitpic[510] <= 4'b1111;
        r_rabbitpic[511] <= 4'b0000;
        r_rabbitpic[512] <= 4'b1111;
        r_rabbitpic[513] <= 4'b1111;
        r_rabbitpic[514] <= 4'b0000;
        r_rabbitpic[515] <= 4'b0000;
        r_rabbitpic[516] <= 4'b1111;
        r_rabbitpic[517] <= 4'b1111;
        r_rabbitpic[518] <= 4'b0000;
        r_rabbitpic[519] <= 4'b0000;
        r_rabbitpic[520] <= 4'b1111;
        r_rabbitpic[521] <= 4'b1111;
        r_rabbitpic[522] <= 4'b0000;
        r_rabbitpic[523] <= 4'b1111;
        r_rabbitpic[524] <= 4'b1111;
        r_rabbitpic[525] <= 4'b1111;
        r_rabbitpic[526] <= 4'b1111;
        r_rabbitpic[527] <= 4'b1111;
        r_rabbitpic[528] <= 4'b1111;
        r_rabbitpic[529] <= 4'b1111;
        r_rabbitpic[530] <= 4'b1111;
        r_rabbitpic[531] <= 4'b1111;
        r_rabbitpic[532] <= 4'b1111;
        r_rabbitpic[533] <= 4'b1111;
        r_rabbitpic[534] <= 4'b1111;
        r_rabbitpic[535] <= 4'b1111;
        r_rabbitpic[536] <= 4'b1111;
        r_rabbitpic[537] <= 4'b1111;
        r_rabbitpic[538] <= 4'b1111;
        r_rabbitpic[539] <= 4'b1111;
        r_rabbitpic[540] <= 4'b1111;
        r_rabbitpic[541] <= 4'b1111;
        r_rabbitpic[542] <= 4'b1111;
        r_rabbitpic[543] <= 4'b1111;
        r_rabbitpic[544] <= 4'b1111;
        r_rabbitpic[545] <= 4'b1111;
        r_rabbitpic[546] <= 4'b1111;
        r_rabbitpic[547] <= 4'b1111;
        r_rabbitpic[548] <= 4'b1111;
        r_rabbitpic[549] <= 4'b1111;
        r_rabbitpic[550] <= 4'b1111;
        r_rabbitpic[551] <= 4'b1111;
        r_rabbitpic[552] <= 4'b1111;
        r_rabbitpic[553] <= 4'b1111;
        r_rabbitpic[554] <= 4'b1111;
        r_rabbitpic[555] <= 4'b1111;
        r_rabbitpic[556] <= 4'b1111;
        r_rabbitpic[557] <= 4'b1111;
        r_rabbitpic[558] <= 4'b1111;
        r_rabbitpic[559] <= 4'b1111;
        r_rabbitpic[560] <= 4'b1111;
        r_rabbitpic[561] <= 4'b1111;
        r_rabbitpic[562] <= 4'b1111;
        r_rabbitpic[563] <= 4'b1111;
        r_rabbitpic[564] <= 4'b1111;
        r_rabbitpic[565] <= 4'b1111;
        r_rabbitpic[566] <= 4'b0000;
        r_rabbitpic[567] <= 4'b1111;
        r_rabbitpic[568] <= 4'b1111;
        r_rabbitpic[569] <= 4'b1111;
        r_rabbitpic[570] <= 4'b0000;
        r_rabbitpic[571] <= 4'b0000;
        r_rabbitpic[572] <= 4'b0000;
        r_rabbitpic[573] <= 4'b0000;
        r_rabbitpic[574] <= 4'b1111;
        r_rabbitpic[575] <= 4'b1111;
        r_rabbitpic[576] <= 4'b1111;
        r_rabbitpic[577] <= 4'b0000;
        r_rabbitpic[578] <= 4'b1111;
        r_rabbitpic[579] <= 4'b1111;
        r_rabbitpic[580] <= 4'b1111;
        r_rabbitpic[581] <= 4'b1111;
        r_rabbitpic[582] <= 4'b1111;
        r_rabbitpic[583] <= 4'b1111;
        r_rabbitpic[584] <= 4'b1111;
        r_rabbitpic[585] <= 4'b1111;
        r_rabbitpic[586] <= 4'b1111;
        r_rabbitpic[587] <= 4'b1111;
        r_rabbitpic[588] <= 4'b1111;
        r_rabbitpic[589] <= 4'b1111;
        r_rabbitpic[590] <= 4'b1111;
        r_rabbitpic[591] <= 4'b1111;
        r_rabbitpic[592] <= 4'b1111;
        r_rabbitpic[593] <= 4'b1111;
        r_rabbitpic[594] <= 4'b1111;
        r_rabbitpic[595] <= 4'b1111;
        r_rabbitpic[596] <= 4'b1111;
        r_rabbitpic[597] <= 4'b1111;
        r_rabbitpic[598] <= 4'b1111;
        r_rabbitpic[599] <= 4'b1111;
        r_rabbitpic[600] <= 4'b1111;
        r_rabbitpic[601] <= 4'b1111;
        r_rabbitpic[602] <= 4'b1111;
        r_rabbitpic[603] <= 4'b1111;
        r_rabbitpic[604] <= 4'b1111;
        r_rabbitpic[605] <= 4'b1111;
        r_rabbitpic[606] <= 4'b1111;
        r_rabbitpic[607] <= 4'b1111;
        r_rabbitpic[608] <= 4'b1111;
        r_rabbitpic[609] <= 4'b1111;
        r_rabbitpic[610] <= 4'b1111;
        r_rabbitpic[611] <= 4'b1111;
        r_rabbitpic[612] <= 4'b1111;
        r_rabbitpic[613] <= 4'b1111;
        r_rabbitpic[614] <= 4'b1111;
        r_rabbitpic[615] <= 4'b1111;
        r_rabbitpic[616] <= 4'b1111;
        r_rabbitpic[617] <= 4'b1111;
        r_rabbitpic[618] <= 4'b1111;
        r_rabbitpic[619] <= 4'b1111;
        r_rabbitpic[620] <= 4'b1111;
        r_rabbitpic[621] <= 4'b1111;
        r_rabbitpic[622] <= 4'b1111;
        r_rabbitpic[623] <= 4'b1111;
        r_rabbitpic[624] <= 4'b1111;
        r_rabbitpic[625] <= 4'b0000;
        r_rabbitpic[626] <= 4'b0000;
        r_rabbitpic[627] <= 4'b0000;
        r_rabbitpic[628] <= 4'b0000;
        r_rabbitpic[629] <= 4'b1111;
        r_rabbitpic[630] <= 4'b1111;
        r_rabbitpic[631] <= 4'b0000;
        r_rabbitpic[632] <= 4'b1111;
        r_rabbitpic[633] <= 4'b1111;
        r_rabbitpic[634] <= 4'b1111;
        r_rabbitpic[635] <= 4'b1111;
        r_rabbitpic[636] <= 4'b1111;
        r_rabbitpic[637] <= 4'b1111;
        r_rabbitpic[638] <= 4'b1111;
        r_rabbitpic[639] <= 4'b1111;
        r_rabbitpic[640] <= 4'b1111;
        r_rabbitpic[641] <= 4'b1111;
        r_rabbitpic[642] <= 4'b1111;
        r_rabbitpic[643] <= 4'b1111;
        r_rabbitpic[644] <= 4'b1111;
        r_rabbitpic[645] <= 4'b1111;
        r_rabbitpic[646] <= 4'b1111;
        r_rabbitpic[647] <= 4'b1111;
        r_rabbitpic[648] <= 4'b1111;
        r_rabbitpic[649] <= 4'b1111;
        r_rabbitpic[650] <= 4'b1111;
        r_rabbitpic[651] <= 4'b1111;
        r_rabbitpic[652] <= 4'b1111;
        r_rabbitpic[653] <= 4'b1111;
        r_rabbitpic[654] <= 4'b1111;
        r_rabbitpic[655] <= 4'b1111;
        r_rabbitpic[656] <= 4'b1111;
        r_rabbitpic[657] <= 4'b1111;
        r_rabbitpic[658] <= 4'b1111;
        r_rabbitpic[659] <= 4'b1111;
        r_rabbitpic[660] <= 4'b1111;
        r_rabbitpic[661] <= 4'b1111;
        r_rabbitpic[662] <= 4'b1111;
        r_rabbitpic[663] <= 4'b1111;
        r_rabbitpic[664] <= 4'b1111;
        r_rabbitpic[665] <= 4'b1111;
        r_rabbitpic[666] <= 4'b1111;
        r_rabbitpic[667] <= 4'b1111;
        r_rabbitpic[668] <= 4'b1111;
        r_rabbitpic[669] <= 4'b1111;
        r_rabbitpic[670] <= 4'b1111;
        r_rabbitpic[671] <= 4'b1111;
        r_rabbitpic[672] <= 4'b1111;
        r_rabbitpic[673] <= 4'b1111;
        r_rabbitpic[674] <= 4'b1111;
        r_rabbitpic[675] <= 4'b1111;
        r_rabbitpic[676] <= 4'b1111;
        r_rabbitpic[677] <= 4'b0000;
        r_rabbitpic[678] <= 4'b1111;
        r_rabbitpic[679] <= 4'b1111;
        r_rabbitpic[680] <= 4'b0000;
        r_rabbitpic[681] <= 4'b0000;
        r_rabbitpic[682] <= 4'b0000;
        r_rabbitpic[683] <= 4'b0000;
        r_rabbitpic[684] <= 4'b1111;
        r_rabbitpic[685] <= 4'b1111;
        r_rabbitpic[686] <= 4'b0000;
        r_rabbitpic[687] <= 4'b1111;
        r_rabbitpic[688] <= 4'b1111;
        r_rabbitpic[689] <= 4'b1111;
        r_rabbitpic[690] <= 4'b1111;
        r_rabbitpic[691] <= 4'b1111;
        r_rabbitpic[692] <= 4'b1111;
        r_rabbitpic[693] <= 4'b1111;
        r_rabbitpic[694] <= 4'b1111;
        r_rabbitpic[695] <= 4'b1111;
        r_rabbitpic[696] <= 4'b1111;
        r_rabbitpic[697] <= 4'b1111;
        r_rabbitpic[698] <= 4'b1111;
        r_rabbitpic[699] <= 4'b1111;
        r_rabbitpic[700] <= 4'b1111;
        r_rabbitpic[701] <= 4'b1111;
        r_rabbitpic[702] <= 4'b1111;
        r_rabbitpic[703] <= 4'b1111;
        r_rabbitpic[704] <= 4'b1111;
        r_rabbitpic[705] <= 4'b1111;
        r_rabbitpic[706] <= 4'b1111;
        r_rabbitpic[707] <= 4'b1111;
        r_rabbitpic[708] <= 4'b1111;
        r_rabbitpic[709] <= 4'b1111;
        r_rabbitpic[710] <= 4'b1111;
        r_rabbitpic[711] <= 4'b1111;
        r_rabbitpic[712] <= 4'b1111;
        r_rabbitpic[713] <= 4'b1111;
        r_rabbitpic[714] <= 4'b1111;
        r_rabbitpic[715] <= 4'b1111;
        r_rabbitpic[716] <= 4'b1111;
        r_rabbitpic[717] <= 4'b1111;
        r_rabbitpic[718] <= 4'b1111;
        r_rabbitpic[719] <= 4'b1111;
        r_rabbitpic[720] <= 4'b1111;
        r_rabbitpic[721] <= 4'b1111;
        r_rabbitpic[722] <= 4'b1111;
        r_rabbitpic[723] <= 4'b1111;
        r_rabbitpic[724] <= 4'b1111;
        r_rabbitpic[725] <= 4'b1111;
        r_rabbitpic[726] <= 4'b1111;
        r_rabbitpic[727] <= 4'b1111;
        r_rabbitpic[728] <= 4'b1111;
        r_rabbitpic[729] <= 4'b1111;
        r_rabbitpic[730] <= 4'b1111;
        r_rabbitpic[731] <= 4'b1111;
        r_rabbitpic[732] <= 4'b0000;
        r_rabbitpic[733] <= 4'b1111;
        r_rabbitpic[734] <= 4'b1111;
        r_rabbitpic[735] <= 4'b1111;
        r_rabbitpic[736] <= 4'b0000;
        r_rabbitpic[737] <= 4'b0000;
        r_rabbitpic[738] <= 4'b1111;
        r_rabbitpic[739] <= 4'b1111;
        r_rabbitpic[740] <= 4'b1111;
        r_rabbitpic[741] <= 4'b0000;
        r_rabbitpic[742] <= 4'b1111;
        r_rabbitpic[743] <= 4'b1111;
        r_rabbitpic[744] <= 4'b1111;
        r_rabbitpic[745] <= 4'b1111;
        r_rabbitpic[746] <= 4'b1111;
        r_rabbitpic[747] <= 4'b1111;
        r_rabbitpic[748] <= 4'b1111;
        r_rabbitpic[749] <= 4'b1111;
        r_rabbitpic[750] <= 4'b1111;
        r_rabbitpic[751] <= 4'b1111;
        r_rabbitpic[752] <= 4'b1111;
        r_rabbitpic[753] <= 4'b1111;
        r_rabbitpic[754] <= 4'b1111;
        r_rabbitpic[755] <= 4'b1111;
        r_rabbitpic[756] <= 4'b1111;
        r_rabbitpic[757] <= 4'b1111;
        r_rabbitpic[758] <= 4'b1111;
        r_rabbitpic[759] <= 4'b1111;
        r_rabbitpic[760] <= 4'b1111;
        r_rabbitpic[761] <= 4'b1111;
        r_rabbitpic[762] <= 4'b1111;
        r_rabbitpic[763] <= 4'b1111;
        r_rabbitpic[764] <= 4'b1111;
        r_rabbitpic[765] <= 4'b1111;
        r_rabbitpic[766] <= 4'b1111;
        r_rabbitpic[767] <= 4'b1111;
        r_rabbitpic[768] <= 4'b1111;
        r_rabbitpic[769] <= 4'b1111;
        r_rabbitpic[770] <= 4'b1111;
        r_rabbitpic[771] <= 4'b1111;
        r_rabbitpic[772] <= 4'b1111;
        r_rabbitpic[773] <= 4'b1111;
        r_rabbitpic[774] <= 4'b1111;
        r_rabbitpic[775] <= 4'b1111;
        r_rabbitpic[776] <= 4'b1111;
        r_rabbitpic[777] <= 4'b1111;
        r_rabbitpic[778] <= 4'b1111;
        r_rabbitpic[779] <= 4'b1111;
        r_rabbitpic[780] <= 4'b1111;
        r_rabbitpic[781] <= 4'b1111;
        r_rabbitpic[782] <= 4'b1111;
        r_rabbitpic[783] <= 4'b1111;
        r_rabbitpic[784] <= 4'b1111;
        r_rabbitpic[785] <= 4'b1111;
        r_rabbitpic[786] <= 4'b1111;
        r_rabbitpic[787] <= 4'b1111;
        r_rabbitpic[788] <= 4'b0000;
        r_rabbitpic[789] <= 4'b1111;
        r_rabbitpic[790] <= 4'b1111;
        r_rabbitpic[791] <= 4'b0000;
        r_rabbitpic[792] <= 4'b0000;
        r_rabbitpic[793] <= 4'b1111;
        r_rabbitpic[794] <= 4'b1111;
        r_rabbitpic[795] <= 4'b0000;
        r_rabbitpic[796] <= 4'b1111;
        r_rabbitpic[797] <= 4'b1111;
        r_rabbitpic[798] <= 4'b1111;
        r_rabbitpic[799] <= 4'b1111;
        r_rabbitpic[800] <= 4'b1111;
        r_rabbitpic[801] <= 4'b1111;
        r_rabbitpic[802] <= 4'b1111;
        r_rabbitpic[803] <= 4'b1111;
        r_rabbitpic[804] <= 4'b1111;
        r_rabbitpic[805] <= 4'b1111;
        r_rabbitpic[806] <= 4'b1111;
        r_rabbitpic[807] <= 4'b1111;
        r_rabbitpic[808] <= 4'b1111;
        r_rabbitpic[809] <= 4'b1111;
        r_rabbitpic[810] <= 4'b1111;
        r_rabbitpic[811] <= 4'b1111;
        r_rabbitpic[812] <= 4'b1111;
        r_rabbitpic[813] <= 4'b1111;
        r_rabbitpic[814] <= 4'b1111;
        r_rabbitpic[815] <= 4'b1111;
        r_rabbitpic[816] <= 4'b1111;
        r_rabbitpic[817] <= 4'b1111;
        r_rabbitpic[818] <= 4'b1111;
        r_rabbitpic[819] <= 4'b1111;
        r_rabbitpic[820] <= 4'b1111;
        r_rabbitpic[821] <= 4'b1111;
        r_rabbitpic[822] <= 4'b1111;
        r_rabbitpic[823] <= 4'b1111;
        r_rabbitpic[824] <= 4'b1111;
        r_rabbitpic[825] <= 4'b1111;
        r_rabbitpic[826] <= 4'b1111;
        r_rabbitpic[827] <= 4'b1111;
        r_rabbitpic[828] <= 4'b1111;
        r_rabbitpic[829] <= 4'b1111;
        r_rabbitpic[830] <= 4'b1111;
        r_rabbitpic[831] <= 4'b1111;
        r_rabbitpic[832] <= 4'b1111;
        r_rabbitpic[833] <= 4'b1111;
        r_rabbitpic[834] <= 4'b1111;
        r_rabbitpic[835] <= 4'b1111;
        r_rabbitpic[836] <= 4'b1111;
        r_rabbitpic[837] <= 4'b1111;
        r_rabbitpic[838] <= 4'b1111;
        r_rabbitpic[839] <= 4'b1111;
        r_rabbitpic[840] <= 4'b1111;
        r_rabbitpic[841] <= 4'b1111;
        r_rabbitpic[842] <= 4'b1111;
        r_rabbitpic[843] <= 4'b0000;
        r_rabbitpic[844] <= 4'b1111;
        r_rabbitpic[845] <= 4'b1111;
        r_rabbitpic[846] <= 4'b0000;
        r_rabbitpic[847] <= 4'b0000;
        r_rabbitpic[848] <= 4'b1111;
        r_rabbitpic[849] <= 4'b1111;
        r_rabbitpic[850] <= 4'b0000;
        r_rabbitpic[851] <= 4'b1111;
        r_rabbitpic[852] <= 4'b1111;
        r_rabbitpic[853] <= 4'b1111;
        r_rabbitpic[854] <= 4'b1111;
        r_rabbitpic[855] <= 4'b1111;
        r_rabbitpic[856] <= 4'b1111;
        r_rabbitpic[857] <= 4'b1111;
        r_rabbitpic[858] <= 4'b1111;
        r_rabbitpic[859] <= 4'b1111;
        r_rabbitpic[860] <= 4'b1111;
        r_rabbitpic[861] <= 4'b1111;
        r_rabbitpic[862] <= 4'b1111;
        r_rabbitpic[863] <= 4'b1111;
        r_rabbitpic[864] <= 4'b1111;
        r_rabbitpic[865] <= 4'b1111;
        r_rabbitpic[866] <= 4'b1111;
        r_rabbitpic[867] <= 4'b1111;
        r_rabbitpic[868] <= 4'b1111;
        r_rabbitpic[869] <= 4'b1111;
        r_rabbitpic[870] <= 4'b1111;
        r_rabbitpic[871] <= 4'b1111;
        r_rabbitpic[872] <= 4'b1111;
        r_rabbitpic[873] <= 4'b1111;
        r_rabbitpic[874] <= 4'b1111;
        r_rabbitpic[875] <= 4'b1111;
        r_rabbitpic[876] <= 4'b1111;
        r_rabbitpic[877] <= 4'b1111;
        r_rabbitpic[878] <= 4'b1111;
        r_rabbitpic[879] <= 4'b1111;
        r_rabbitpic[880] <= 4'b1111;
        r_rabbitpic[881] <= 4'b1111;
        r_rabbitpic[882] <= 4'b1111;
        r_rabbitpic[883] <= 4'b1111;
        r_rabbitpic[884] <= 4'b1111;
        r_rabbitpic[885] <= 4'b1111;
        r_rabbitpic[886] <= 4'b1111;
        r_rabbitpic[887] <= 4'b1111;
        r_rabbitpic[888] <= 4'b1111;
        r_rabbitpic[889] <= 4'b1111;
        r_rabbitpic[890] <= 4'b1111;
        r_rabbitpic[891] <= 4'b1111;
        r_rabbitpic[892] <= 4'b1111;
        r_rabbitpic[893] <= 4'b1111;
        r_rabbitpic[894] <= 4'b1111;
        r_rabbitpic[895] <= 4'b1111;
        r_rabbitpic[896] <= 4'b1111;
        r_rabbitpic[897] <= 4'b1111;
        r_rabbitpic[898] <= 4'b1111;
        r_rabbitpic[899] <= 4'b0000;
        r_rabbitpic[900] <= 4'b0000;
        r_rabbitpic[901] <= 4'b0000;
        r_rabbitpic[902] <= 4'b0000;
        r_rabbitpic[903] <= 4'b0000;
        r_rabbitpic[904] <= 4'b0000;
        r_rabbitpic[905] <= 4'b1111;
        r_rabbitpic[906] <= 4'b1111;
        r_rabbitpic[907] <= 4'b1111;
        r_rabbitpic[908] <= 4'b1111;
        r_rabbitpic[909] <= 4'b1111;
        r_rabbitpic[910] <= 4'b1111;
        r_rabbitpic[911] <= 4'b1111;
        r_rabbitpic[912] <= 4'b1111;
        r_rabbitpic[913] <= 4'b1111;
        r_rabbitpic[914] <= 4'b1111;
        r_rabbitpic[915] <= 4'b1111;
        r_rabbitpic[916] <= 4'b1111;
        r_rabbitpic[917] <= 4'b1111;
        r_rabbitpic[918] <= 4'b1111;
        r_rabbitpic[919] <= 4'b1111;
        r_rabbitpic[920] <= 4'b1111;
        r_rabbitpic[921] <= 4'b1111;
        r_rabbitpic[922] <= 4'b1111;
        r_rabbitpic[923] <= 4'b1111;
        r_rabbitpic[924] <= 4'b1111;
        r_rabbitpic[925] <= 4'b1111;
        r_rabbitpic[926] <= 4'b1111;
        r_rabbitpic[927] <= 4'b1111;
        r_rabbitpic[928] <= 4'b1111;
        r_rabbitpic[929] <= 4'b1111;
        r_rabbitpic[930] <= 4'b1111;
        r_rabbitpic[931] <= 4'b1111;
        r_rabbitpic[932] <= 4'b1111;
        r_rabbitpic[933] <= 4'b1111;
        r_rabbitpic[934] <= 4'b1111;
        r_rabbitpic[935] <= 4'b1111;
        r_rabbitpic[936] <= 4'b1111;
        r_rabbitpic[937] <= 4'b1111;
        r_rabbitpic[938] <= 4'b1111;
        r_rabbitpic[939] <= 4'b1111;
        r_rabbitpic[940] <= 4'b1111;
        r_rabbitpic[941] <= 4'b1111;
        r_rabbitpic[942] <= 4'b1111;
        r_rabbitpic[943] <= 4'b1111;
        r_rabbitpic[944] <= 4'b1111;
        r_rabbitpic[945] <= 4'b1111;
        r_rabbitpic[946] <= 4'b1111;
        r_rabbitpic[947] <= 4'b1111;
        r_rabbitpic[948] <= 4'b1111;
        r_rabbitpic[949] <= 4'b1111;
        r_rabbitpic[950] <= 4'b1111;
        r_rabbitpic[951] <= 4'b1111;
        r_rabbitpic[952] <= 4'b1111;
        r_rabbitpic[953] <= 4'b1111;
        r_rabbitpic[954] <= 4'b0000;
        r_rabbitpic[955] <= 4'b1111;
        r_rabbitpic[956] <= 4'b1111;
        r_rabbitpic[957] <= 4'b1111;
        r_rabbitpic[958] <= 4'b1111;
        r_rabbitpic[959] <= 4'b0000;
        r_rabbitpic[960] <= 4'b1111;
        r_rabbitpic[961] <= 4'b1111;
        r_rabbitpic[962] <= 4'b1111;
        r_rabbitpic[963] <= 4'b1111;
        r_rabbitpic[964] <= 4'b1111;
        r_rabbitpic[965] <= 4'b1111;
        r_rabbitpic[966] <= 4'b1111;
        r_rabbitpic[967] <= 4'b1111;
        r_rabbitpic[968] <= 4'b1111;
        r_rabbitpic[969] <= 4'b1111;
        r_rabbitpic[970] <= 4'b1111;
        r_rabbitpic[971] <= 4'b1111;
        r_rabbitpic[972] <= 4'b1111;
        r_rabbitpic[973] <= 4'b1111;
        r_rabbitpic[974] <= 4'b1111;
        r_rabbitpic[975] <= 4'b1111;
        r_rabbitpic[976] <= 4'b1111;
        r_rabbitpic[977] <= 4'b1111;
        r_rabbitpic[978] <= 4'b1111;
        r_rabbitpic[979] <= 4'b1111;
        r_rabbitpic[980] <= 4'b1111;
        r_rabbitpic[981] <= 4'b1111;
        r_rabbitpic[982] <= 4'b1111;
        r_rabbitpic[983] <= 4'b1111;
        r_rabbitpic[984] <= 4'b1111;
        r_rabbitpic[985] <= 4'b1111;
        r_rabbitpic[986] <= 4'b1111;
        r_rabbitpic[987] <= 4'b1111;
        r_rabbitpic[988] <= 4'b1111;
        r_rabbitpic[989] <= 4'b1111;
        r_rabbitpic[990] <= 4'b1111;
        r_rabbitpic[991] <= 4'b1111;
        r_rabbitpic[992] <= 4'b1111;
        r_rabbitpic[993] <= 4'b1111;
        r_rabbitpic[994] <= 4'b1111;
        r_rabbitpic[995] <= 4'b1111;
        r_rabbitpic[996] <= 4'b1111;
        r_rabbitpic[997] <= 4'b1111;
        r_rabbitpic[998] <= 4'b1111;
        r_rabbitpic[999] <= 4'b1111;
        r_rabbitpic[1000] <= 4'b1111;
        r_rabbitpic[1001] <= 4'b1111;
        r_rabbitpic[1002] <= 4'b1111;
        r_rabbitpic[1003] <= 4'b1111;
        r_rabbitpic[1004] <= 4'b1111;
        r_rabbitpic[1005] <= 4'b1111;
        r_rabbitpic[1006] <= 4'b1111;
        r_rabbitpic[1007] <= 4'b1111;
        r_rabbitpic[1008] <= 4'b0000;
        r_rabbitpic[1009] <= 4'b1111;
        r_rabbitpic[1010] <= 4'b1111;
        r_rabbitpic[1011] <= 4'b1111;
        r_rabbitpic[1012] <= 4'b1111;
        r_rabbitpic[1013] <= 4'b1111;
        r_rabbitpic[1014] <= 4'b1111;
        r_rabbitpic[1015] <= 4'b0000;
        r_rabbitpic[1016] <= 4'b1111;
        r_rabbitpic[1017] <= 4'b1111;
        r_rabbitpic[1018] <= 4'b1111;
        r_rabbitpic[1019] <= 4'b1111;
        r_rabbitpic[1020] <= 4'b1111;
        r_rabbitpic[1021] <= 4'b1111;
        r_rabbitpic[1022] <= 4'b1111;
        r_rabbitpic[1023] <= 4'b1111;
        r_rabbitpic[1024] <= 4'b1111;
        r_rabbitpic[1025] <= 4'b1111;
        r_rabbitpic[1026] <= 4'b1111;
        r_rabbitpic[1027] <= 4'b1111;
        r_rabbitpic[1028] <= 4'b1111;
        r_rabbitpic[1029] <= 4'b1111;
        r_rabbitpic[1030] <= 4'b1111;
        r_rabbitpic[1031] <= 4'b1111;
        r_rabbitpic[1032] <= 4'b1111;
        r_rabbitpic[1033] <= 4'b1111;
        r_rabbitpic[1034] <= 4'b1111;
        r_rabbitpic[1035] <= 4'b1111;
        r_rabbitpic[1036] <= 4'b1111;
        r_rabbitpic[1037] <= 4'b1111;
        r_rabbitpic[1038] <= 4'b1111;
        r_rabbitpic[1039] <= 4'b1111;
        r_rabbitpic[1040] <= 4'b1111;
        r_rabbitpic[1041] <= 4'b1111;
        r_rabbitpic[1042] <= 4'b1111;
        r_rabbitpic[1043] <= 4'b1111;
        r_rabbitpic[1044] <= 4'b1111;
        r_rabbitpic[1045] <= 4'b1111;
        r_rabbitpic[1046] <= 4'b1111;
        r_rabbitpic[1047] <= 4'b1111;
        r_rabbitpic[1048] <= 4'b1111;
        r_rabbitpic[1049] <= 4'b1111;
        r_rabbitpic[1050] <= 4'b1111;
        r_rabbitpic[1051] <= 4'b1111;
        r_rabbitpic[1052] <= 4'b1111;
        r_rabbitpic[1053] <= 4'b1111;
        r_rabbitpic[1054] <= 4'b1111;
        r_rabbitpic[1055] <= 4'b1111;
        r_rabbitpic[1056] <= 4'b1111;
        r_rabbitpic[1057] <= 4'b1111;
        r_rabbitpic[1058] <= 4'b1111;
        r_rabbitpic[1059] <= 4'b1111;
        r_rabbitpic[1060] <= 4'b1111;
        r_rabbitpic[1061] <= 4'b1111;
        r_rabbitpic[1062] <= 4'b1111;
        r_rabbitpic[1063] <= 4'b0000;
        r_rabbitpic[1064] <= 4'b0000;
        r_rabbitpic[1065] <= 4'b0000;
        r_rabbitpic[1066] <= 4'b1111;
        r_rabbitpic[1067] <= 4'b1111;
        r_rabbitpic[1068] <= 4'b1111;
        r_rabbitpic[1069] <= 4'b0000;
        r_rabbitpic[1070] <= 4'b0000;
        r_rabbitpic[1071] <= 4'b0000;
        r_rabbitpic[1072] <= 4'b1111;
        r_rabbitpic[1073] <= 4'b1111;
        r_rabbitpic[1074] <= 4'b1111;
        r_rabbitpic[1075] <= 4'b1111;
        r_rabbitpic[1076] <= 4'b1111;
        r_rabbitpic[1077] <= 4'b1111;
        r_rabbitpic[1078] <= 4'b1111;
        r_rabbitpic[1079] <= 4'b1111;
        r_rabbitpic[1080] <= 4'b1111;
        r_rabbitpic[1081] <= 4'b1111;
        r_rabbitpic[1082] <= 4'b1111;
        r_rabbitpic[1083] <= 4'b1111;
        r_rabbitpic[1084] <= 4'b1111;
        r_rabbitpic[1085] <= 4'b1111;
        r_rabbitpic[1086] <= 4'b1111;
        r_rabbitpic[1087] <= 4'b1111;
        r_rabbitpic[1088] <= 4'b1111;
        r_rabbitpic[1089] <= 4'b1111;
        r_rabbitpic[1090] <= 4'b1111;
        r_rabbitpic[1091] <= 4'b1111;
        r_rabbitpic[1092] <= 4'b1111;
        r_rabbitpic[1093] <= 4'b1111;
        r_rabbitpic[1094] <= 4'b1111;
        r_rabbitpic[1095] <= 4'b1111;
        r_rabbitpic[1096] <= 4'b1111;
        r_rabbitpic[1097] <= 4'b1111;
        r_rabbitpic[1098] <= 4'b1111;
        r_rabbitpic[1099] <= 4'b1111;
        r_rabbitpic[1100] <= 4'b1111;
        r_rabbitpic[1101] <= 4'b1111;
        r_rabbitpic[1102] <= 4'b1111;
        r_rabbitpic[1103] <= 4'b1111;
        r_rabbitpic[1104] <= 4'b1111;
        r_rabbitpic[1105] <= 4'b1111;
        r_rabbitpic[1106] <= 4'b1111;
        r_rabbitpic[1107] <= 4'b1111;
        r_rabbitpic[1108] <= 4'b1111;
        r_rabbitpic[1109] <= 4'b1111;
        r_rabbitpic[1110] <= 4'b1111;
        r_rabbitpic[1111] <= 4'b1111;
        r_rabbitpic[1112] <= 4'b1111;
        r_rabbitpic[1113] <= 4'b1111;
        r_rabbitpic[1114] <= 4'b1111;
        r_rabbitpic[1115] <= 4'b1111;
        r_rabbitpic[1116] <= 4'b1111;
        r_rabbitpic[1117] <= 4'b0000;
        r_rabbitpic[1118] <= 4'b1111;
        r_rabbitpic[1119] <= 4'b0000;
        r_rabbitpic[1120] <= 4'b0000;
        r_rabbitpic[1121] <= 4'b1111;
        r_rabbitpic[1122] <= 4'b1111;
        r_rabbitpic[1123] <= 4'b1111;
        r_rabbitpic[1124] <= 4'b0000;
        r_rabbitpic[1125] <= 4'b1111;
        r_rabbitpic[1126] <= 4'b0000;
        r_rabbitpic[1127] <= 4'b1111;
        r_rabbitpic[1128] <= 4'b1111;
        r_rabbitpic[1129] <= 4'b1111;
        r_rabbitpic[1130] <= 4'b1111;
        r_rabbitpic[1131] <= 4'b1111;
        r_rabbitpic[1132] <= 4'b1111;
        r_rabbitpic[1133] <= 4'b1111;
        r_rabbitpic[1134] <= 4'b1111;
        r_rabbitpic[1135] <= 4'b1111;
        r_rabbitpic[1136] <= 4'b1111;
        r_rabbitpic[1137] <= 4'b1111;
        r_rabbitpic[1138] <= 4'b1111;
        r_rabbitpic[1139] <= 4'b1111;
        r_rabbitpic[1140] <= 4'b1111;
        r_rabbitpic[1141] <= 4'b1111;
        r_rabbitpic[1142] <= 4'b1111;
        r_rabbitpic[1143] <= 4'b1111;
        r_rabbitpic[1144] <= 4'b1111;
        r_rabbitpic[1145] <= 4'b1111;
        r_rabbitpic[1146] <= 4'b1111;
        r_rabbitpic[1147] <= 4'b1111;
        r_rabbitpic[1148] <= 4'b1111;
        r_rabbitpic[1149] <= 4'b1111;
        r_rabbitpic[1150] <= 4'b1111;
        r_rabbitpic[1151] <= 4'b1111;
        r_rabbitpic[1152] <= 4'b1111;
        r_rabbitpic[1153] <= 4'b1111;
        r_rabbitpic[1154] <= 4'b1111;
        r_rabbitpic[1155] <= 4'b1111;
        r_rabbitpic[1156] <= 4'b1111;
        r_rabbitpic[1157] <= 4'b1111;
        r_rabbitpic[1158] <= 4'b1111;
        r_rabbitpic[1159] <= 4'b1111;
        r_rabbitpic[1160] <= 4'b1111;
        r_rabbitpic[1161] <= 4'b1111;
        r_rabbitpic[1162] <= 4'b1111;
        r_rabbitpic[1163] <= 4'b1111;
        r_rabbitpic[1164] <= 4'b1111;
        r_rabbitpic[1165] <= 4'b1111;
        r_rabbitpic[1166] <= 4'b1111;
        r_rabbitpic[1167] <= 4'b1111;
        r_rabbitpic[1168] <= 4'b1111;
        r_rabbitpic[1169] <= 4'b1111;
        r_rabbitpic[1170] <= 4'b1111;
        r_rabbitpic[1171] <= 4'b1111;
        r_rabbitpic[1172] <= 4'b0000;
        r_rabbitpic[1173] <= 4'b1111;
        r_rabbitpic[1174] <= 4'b1111;
        r_rabbitpic[1175] <= 4'b1111;
        r_rabbitpic[1176] <= 4'b1111;
        r_rabbitpic[1177] <= 4'b1111;
        r_rabbitpic[1178] <= 4'b1111;
        r_rabbitpic[1179] <= 4'b1111;
        r_rabbitpic[1180] <= 4'b1111;
        r_rabbitpic[1181] <= 4'b1111;
        r_rabbitpic[1182] <= 4'b0000;
        r_rabbitpic[1183] <= 4'b1111;
        r_rabbitpic[1184] <= 4'b1111;
        r_rabbitpic[1185] <= 4'b1111;
        r_rabbitpic[1186] <= 4'b1111;
        r_rabbitpic[1187] <= 4'b1111;
        r_rabbitpic[1188] <= 4'b1111;
        r_rabbitpic[1189] <= 4'b1111;
        r_rabbitpic[1190] <= 4'b1111;
        r_rabbitpic[1191] <= 4'b1111;
        r_rabbitpic[1192] <= 4'b1111;
        r_rabbitpic[1193] <= 4'b1111;
        r_rabbitpic[1194] <= 4'b1111;
        r_rabbitpic[1195] <= 4'b1111;
        r_rabbitpic[1196] <= 4'b1111;
        r_rabbitpic[1197] <= 4'b1111;
        r_rabbitpic[1198] <= 4'b1111;
        r_rabbitpic[1199] <= 4'b1111;
        r_rabbitpic[1200] <= 4'b1111;
        r_rabbitpic[1201] <= 4'b1111;
        r_rabbitpic[1202] <= 4'b1111;
        r_rabbitpic[1203] <= 4'b1111;
        r_rabbitpic[1204] <= 4'b1111;
        r_rabbitpic[1205] <= 4'b1111;
        r_rabbitpic[1206] <= 4'b1111;
        r_rabbitpic[1207] <= 4'b1111;
        r_rabbitpic[1208] <= 4'b1111;
        r_rabbitpic[1209] <= 4'b1111;
        r_rabbitpic[1210] <= 4'b1111;
        r_rabbitpic[1211] <= 4'b1111;
        r_rabbitpic[1212] <= 4'b1111;
        r_rabbitpic[1213] <= 4'b1111;
        r_rabbitpic[1214] <= 4'b1111;
        r_rabbitpic[1215] <= 4'b1111;
        r_rabbitpic[1216] <= 4'b1111;
        r_rabbitpic[1217] <= 4'b1111;
        r_rabbitpic[1218] <= 4'b1111;
        r_rabbitpic[1219] <= 4'b1111;
        r_rabbitpic[1220] <= 4'b1111;
        r_rabbitpic[1221] <= 4'b1111;
        r_rabbitpic[1222] <= 4'b1111;
        r_rabbitpic[1223] <= 4'b1111;
        r_rabbitpic[1224] <= 4'b1111;
        r_rabbitpic[1225] <= 4'b1111;
        r_rabbitpic[1226] <= 4'b1111;
        r_rabbitpic[1227] <= 4'b0000;
        r_rabbitpic[1228] <= 4'b1111;
        r_rabbitpic[1229] <= 4'b1111;
        r_rabbitpic[1230] <= 4'b1111;
        r_rabbitpic[1231] <= 4'b1111;
        r_rabbitpic[1232] <= 4'b1111;
        r_rabbitpic[1233] <= 4'b1111;
        r_rabbitpic[1234] <= 4'b1111;
        r_rabbitpic[1235] <= 4'b1111;
        r_rabbitpic[1236] <= 4'b1111;
        r_rabbitpic[1237] <= 4'b0000;
        r_rabbitpic[1238] <= 4'b1111;
        r_rabbitpic[1239] <= 4'b1111;
        r_rabbitpic[1240] <= 4'b1111;
        r_rabbitpic[1241] <= 4'b1111;
        r_rabbitpic[1242] <= 4'b1111;
        r_rabbitpic[1243] <= 4'b1111;
        r_rabbitpic[1244] <= 4'b1111;
        r_rabbitpic[1245] <= 4'b1111;
        r_rabbitpic[1246] <= 4'b1111;
        r_rabbitpic[1247] <= 4'b1111;
        r_rabbitpic[1248] <= 4'b1111;
        r_rabbitpic[1249] <= 4'b1111;
        r_rabbitpic[1250] <= 4'b1111;
        r_rabbitpic[1251] <= 4'b1111;
        r_rabbitpic[1252] <= 4'b1111;
        r_rabbitpic[1253] <= 4'b1111;
        r_rabbitpic[1254] <= 4'b1111;
        r_rabbitpic[1255] <= 4'b1111;
        r_rabbitpic[1256] <= 4'b1111;
        r_rabbitpic[1257] <= 4'b1111;
        r_rabbitpic[1258] <= 4'b1111;
        r_rabbitpic[1259] <= 4'b1111;
        r_rabbitpic[1260] <= 4'b1111;
        r_rabbitpic[1261] <= 4'b1111;
        r_rabbitpic[1262] <= 4'b1111;
        r_rabbitpic[1263] <= 4'b1111;
        r_rabbitpic[1264] <= 4'b1111;
        r_rabbitpic[1265] <= 4'b1111;
        r_rabbitpic[1266] <= 4'b1111;
        r_rabbitpic[1267] <= 4'b1111;
        r_rabbitpic[1268] <= 4'b1111;
        r_rabbitpic[1269] <= 4'b1111;
        r_rabbitpic[1270] <= 4'b1111;
        r_rabbitpic[1271] <= 4'b1111;
        r_rabbitpic[1272] <= 4'b1111;
        r_rabbitpic[1273] <= 4'b1111;
        r_rabbitpic[1274] <= 4'b1111;
        r_rabbitpic[1275] <= 4'b1111;
        r_rabbitpic[1276] <= 4'b1111;
        r_rabbitpic[1277] <= 4'b1111;
        r_rabbitpic[1278] <= 4'b1111;
        r_rabbitpic[1279] <= 4'b1111;
        r_rabbitpic[1280] <= 4'b1111;
        r_rabbitpic[1281] <= 4'b0000;
        r_rabbitpic[1282] <= 4'b0000;
        r_rabbitpic[1283] <= 4'b1111;
        r_rabbitpic[1284] <= 4'b1111;
        r_rabbitpic[1285] <= 4'b1111;
        r_rabbitpic[1286] <= 4'b0000;
        r_rabbitpic[1287] <= 4'b0000;
        r_rabbitpic[1288] <= 4'b1111;
        r_rabbitpic[1289] <= 4'b1111;
        r_rabbitpic[1290] <= 4'b1111;
        r_rabbitpic[1291] <= 4'b0000;
        r_rabbitpic[1292] <= 4'b0000;
        r_rabbitpic[1293] <= 4'b1111;
        r_rabbitpic[1294] <= 4'b1111;
        r_rabbitpic[1295] <= 4'b1111;
        r_rabbitpic[1296] <= 4'b1111;
        r_rabbitpic[1297] <= 4'b1111;
        r_rabbitpic[1298] <= 4'b1111;
        r_rabbitpic[1299] <= 4'b1111;
        r_rabbitpic[1300] <= 4'b1111;
        r_rabbitpic[1301] <= 4'b1111;
        r_rabbitpic[1302] <= 4'b1111;
        r_rabbitpic[1303] <= 4'b1111;
        r_rabbitpic[1304] <= 4'b1111;
        r_rabbitpic[1305] <= 4'b1111;
        r_rabbitpic[1306] <= 4'b1111;
        r_rabbitpic[1307] <= 4'b1111;
        r_rabbitpic[1308] <= 4'b1111;
        r_rabbitpic[1309] <= 4'b1111;
        r_rabbitpic[1310] <= 4'b1111;
        r_rabbitpic[1311] <= 4'b1111;
        r_rabbitpic[1312] <= 4'b1111;
        r_rabbitpic[1313] <= 4'b1111;
        r_rabbitpic[1314] <= 4'b1111;
        r_rabbitpic[1315] <= 4'b1111;
        r_rabbitpic[1316] <= 4'b1111;
        r_rabbitpic[1317] <= 4'b1111;
        r_rabbitpic[1318] <= 4'b1111;
        r_rabbitpic[1319] <= 4'b1111;
        r_rabbitpic[1320] <= 4'b1111;
        r_rabbitpic[1321] <= 4'b1111;
        r_rabbitpic[1322] <= 4'b1111;
        r_rabbitpic[1323] <= 4'b1111;
        r_rabbitpic[1324] <= 4'b1111;
        r_rabbitpic[1325] <= 4'b1111;
        r_rabbitpic[1326] <= 4'b1111;
        r_rabbitpic[1327] <= 4'b1111;
        r_rabbitpic[1328] <= 4'b1111;
        r_rabbitpic[1329] <= 4'b1111;
        r_rabbitpic[1330] <= 4'b1111;
        r_rabbitpic[1331] <= 4'b1111;
        r_rabbitpic[1332] <= 4'b1111;
        r_rabbitpic[1333] <= 4'b1111;
        r_rabbitpic[1334] <= 4'b1111;
        r_rabbitpic[1335] <= 4'b1111;
        r_rabbitpic[1336] <= 4'b1111;
        r_rabbitpic[1337] <= 4'b0000;
        r_rabbitpic[1338] <= 4'b1111;
        r_rabbitpic[1339] <= 4'b1111;
        r_rabbitpic[1340] <= 4'b0000;
        r_rabbitpic[1341] <= 4'b0000;
        r_rabbitpic[1342] <= 4'b0000;
        r_rabbitpic[1343] <= 4'b0000;
        r_rabbitpic[1344] <= 4'b1111;
        r_rabbitpic[1345] <= 4'b1111;
        r_rabbitpic[1346] <= 4'b0000;
        r_rabbitpic[1347] <= 4'b0000;
        r_rabbitpic[1348] <= 4'b1111;
        r_rabbitpic[1349] <= 4'b1111;
        r_rabbitpic[1350] <= 4'b1111;
        r_rabbitpic[1351] <= 4'b1111;
        r_rabbitpic[1352] <= 4'b1111;
        r_rabbitpic[1353] <= 4'b1111;
        r_rabbitpic[1354] <= 4'b1111;
        r_rabbitpic[1355] <= 4'b1111;
        r_rabbitpic[1356] <= 4'b1111;
        r_rabbitpic[1357] <= 4'b1111;
        r_rabbitpic[1358] <= 4'b1111;
        r_rabbitpic[1359] <= 4'b1111;
        r_rabbitpic[1360] <= 4'b1111;
        r_rabbitpic[1361] <= 4'b1111;
        r_rabbitpic[1362] <= 4'b1111;
        r_rabbitpic[1363] <= 4'b1111;
        r_rabbitpic[1364] <= 4'b1111;
        r_rabbitpic[1365] <= 4'b1111;
        r_rabbitpic[1366] <= 4'b1111;
        r_rabbitpic[1367] <= 4'b1111;
        r_rabbitpic[1368] <= 4'b1111;
        r_rabbitpic[1369] <= 4'b1111;
        r_rabbitpic[1370] <= 4'b1111;
        r_rabbitpic[1371] <= 4'b1111;
        r_rabbitpic[1372] <= 4'b1111;
        r_rabbitpic[1373] <= 4'b1111;
        r_rabbitpic[1374] <= 4'b1111;
        r_rabbitpic[1375] <= 4'b1111;
        r_rabbitpic[1376] <= 4'b1111;
        r_rabbitpic[1377] <= 4'b1111;
        r_rabbitpic[1378] <= 4'b1111;
        r_rabbitpic[1379] <= 4'b1111;
        r_rabbitpic[1380] <= 4'b1111;
        r_rabbitpic[1381] <= 4'b1111;
        r_rabbitpic[1382] <= 4'b1111;
        r_rabbitpic[1383] <= 4'b1111;
        r_rabbitpic[1384] <= 4'b1111;
        r_rabbitpic[1385] <= 4'b1111;
        r_rabbitpic[1386] <= 4'b1111;
        r_rabbitpic[1387] <= 4'b1111;
        r_rabbitpic[1388] <= 4'b1111;
        r_rabbitpic[1389] <= 4'b1111;
        r_rabbitpic[1390] <= 4'b1111;
        r_rabbitpic[1391] <= 4'b1111;
        r_rabbitpic[1392] <= 4'b1111;
        r_rabbitpic[1393] <= 4'b0000;
        r_rabbitpic[1394] <= 4'b0000;
        r_rabbitpic[1395] <= 4'b1111;
        r_rabbitpic[1396] <= 4'b1111;
        r_rabbitpic[1397] <= 4'b1111;
        r_rabbitpic[1398] <= 4'b1111;
        r_rabbitpic[1399] <= 4'b1111;
        r_rabbitpic[1400] <= 4'b0000;
        r_rabbitpic[1401] <= 4'b1111;
        r_rabbitpic[1402] <= 4'b0000;
        r_rabbitpic[1403] <= 4'b0000;
        r_rabbitpic[1404] <= 4'b1111;
        r_rabbitpic[1405] <= 4'b1111;
        r_rabbitpic[1406] <= 4'b1111;
        r_rabbitpic[1407] <= 4'b1111;
        r_rabbitpic[1408] <= 4'b1111;
        r_rabbitpic[1409] <= 4'b1111;
        r_rabbitpic[1410] <= 4'b1111;
        r_rabbitpic[1411] <= 4'b1111;
        r_rabbitpic[1412] <= 4'b1111;
        r_rabbitpic[1413] <= 4'b1111;
        r_rabbitpic[1414] <= 4'b1111;
        r_rabbitpic[1415] <= 4'b1111;
        r_rabbitpic[1416] <= 4'b1111;
        r_rabbitpic[1417] <= 4'b1111;
        r_rabbitpic[1418] <= 4'b1111;
        r_rabbitpic[1419] <= 4'b1111;
        r_rabbitpic[1420] <= 4'b1111;
        r_rabbitpic[1421] <= 4'b1111;
        r_rabbitpic[1422] <= 4'b1111;
        r_rabbitpic[1423] <= 4'b1111;
        r_rabbitpic[1424] <= 4'b1111;
        r_rabbitpic[1425] <= 4'b1111;
        r_rabbitpic[1426] <= 4'b1111;
        r_rabbitpic[1427] <= 4'b1111;
        r_rabbitpic[1428] <= 4'b1111;
        r_rabbitpic[1429] <= 4'b1111;
        r_rabbitpic[1430] <= 4'b1111;
        r_rabbitpic[1431] <= 4'b1111;
        r_rabbitpic[1432] <= 4'b1111;
        r_rabbitpic[1433] <= 4'b1111;
        r_rabbitpic[1434] <= 4'b1111;
        r_rabbitpic[1435] <= 4'b1111;
        r_rabbitpic[1436] <= 4'b1111;
        r_rabbitpic[1437] <= 4'b1111;
        r_rabbitpic[1438] <= 4'b1111;
        r_rabbitpic[1439] <= 4'b1111;
        r_rabbitpic[1440] <= 4'b1111;
        r_rabbitpic[1441] <= 4'b1111;
        r_rabbitpic[1442] <= 4'b1111;
        r_rabbitpic[1443] <= 4'b1111;
        r_rabbitpic[1444] <= 4'b1111;
        r_rabbitpic[1445] <= 4'b1111;
        r_rabbitpic[1446] <= 4'b1111;
        r_rabbitpic[1447] <= 4'b1111;
        r_rabbitpic[1448] <= 4'b0000;
        r_rabbitpic[1449] <= 4'b1111;
        r_rabbitpic[1450] <= 4'b1111;
        r_rabbitpic[1451] <= 4'b1111;
        r_rabbitpic[1452] <= 4'b1111;
        r_rabbitpic[1453] <= 4'b1111;
        r_rabbitpic[1454] <= 4'b1111;
        r_rabbitpic[1455] <= 4'b1111;
        r_rabbitpic[1456] <= 4'b1111;
        r_rabbitpic[1457] <= 4'b1111;
        r_rabbitpic[1458] <= 4'b1111;
        r_rabbitpic[1459] <= 4'b0000;
        r_rabbitpic[1460] <= 4'b0000;
        r_rabbitpic[1461] <= 4'b1111;
        r_rabbitpic[1462] <= 4'b1111;
        r_rabbitpic[1463] <= 4'b1111;
        r_rabbitpic[1464] <= 4'b1111;
        r_rabbitpic[1465] <= 4'b1111;
        r_rabbitpic[1466] <= 4'b1111;
        r_rabbitpic[1467] <= 4'b1111;
        r_rabbitpic[1468] <= 4'b1111;
        r_rabbitpic[1469] <= 4'b1111;
        r_rabbitpic[1470] <= 4'b1111;
        r_rabbitpic[1471] <= 4'b1111;
        r_rabbitpic[1472] <= 4'b1111;
        r_rabbitpic[1473] <= 4'b1111;
        r_rabbitpic[1474] <= 4'b1111;
        r_rabbitpic[1475] <= 4'b1111;
        r_rabbitpic[1476] <= 4'b1111;
        r_rabbitpic[1477] <= 4'b1111;
        r_rabbitpic[1478] <= 4'b1111;
        r_rabbitpic[1479] <= 4'b1111;
        r_rabbitpic[1480] <= 4'b1111;
        r_rabbitpic[1481] <= 4'b1111;
        r_rabbitpic[1482] <= 4'b1111;
        r_rabbitpic[1483] <= 4'b1111;
        r_rabbitpic[1484] <= 4'b1111;
        r_rabbitpic[1485] <= 4'b1111;
        r_rabbitpic[1486] <= 4'b1111;
        r_rabbitpic[1487] <= 4'b1111;
        r_rabbitpic[1488] <= 4'b1111;
        r_rabbitpic[1489] <= 4'b1111;
        r_rabbitpic[1490] <= 4'b1111;
        r_rabbitpic[1491] <= 4'b1111;
        r_rabbitpic[1492] <= 4'b1111;
        r_rabbitpic[1493] <= 4'b1111;
        r_rabbitpic[1494] <= 4'b1111;
        r_rabbitpic[1495] <= 4'b1111;
        r_rabbitpic[1496] <= 4'b1111;
        r_rabbitpic[1497] <= 4'b1111;
        r_rabbitpic[1498] <= 4'b1111;
        r_rabbitpic[1499] <= 4'b1111;
        r_rabbitpic[1500] <= 4'b1111;
        r_rabbitpic[1501] <= 4'b1111;
        r_rabbitpic[1502] <= 4'b1111;
        r_rabbitpic[1503] <= 4'b0000;
        r_rabbitpic[1504] <= 4'b1111;
        r_rabbitpic[1505] <= 4'b1111;
        r_rabbitpic[1506] <= 4'b1111;
        r_rabbitpic[1507] <= 4'b1111;
        r_rabbitpic[1508] <= 4'b1111;
        r_rabbitpic[1509] <= 4'b1111;
        r_rabbitpic[1510] <= 4'b1111;
        r_rabbitpic[1511] <= 4'b1111;
        r_rabbitpic[1512] <= 4'b1111;
        r_rabbitpic[1513] <= 4'b1111;
        r_rabbitpic[1514] <= 4'b1111;
        r_rabbitpic[1515] <= 4'b1111;
        r_rabbitpic[1516] <= 4'b0000;
        r_rabbitpic[1517] <= 4'b0000;
        r_rabbitpic[1518] <= 4'b0000;
        r_rabbitpic[1519] <= 4'b1111;
        r_rabbitpic[1520] <= 4'b1111;
        r_rabbitpic[1521] <= 4'b1111;
        r_rabbitpic[1522] <= 4'b1111;
        r_rabbitpic[1523] <= 4'b1111;
        r_rabbitpic[1524] <= 4'b1111;
        r_rabbitpic[1525] <= 4'b1111;
        r_rabbitpic[1526] <= 4'b1111;
        r_rabbitpic[1527] <= 4'b1111;
        r_rabbitpic[1528] <= 4'b1111;
        r_rabbitpic[1529] <= 4'b1111;
        r_rabbitpic[1530] <= 4'b1111;
        r_rabbitpic[1531] <= 4'b1111;
        r_rabbitpic[1532] <= 4'b1111;
        r_rabbitpic[1533] <= 4'b1111;
        r_rabbitpic[1534] <= 4'b1111;
        r_rabbitpic[1535] <= 4'b1111;
        r_rabbitpic[1536] <= 4'b1111;
        r_rabbitpic[1537] <= 4'b1111;
        r_rabbitpic[1538] <= 4'b1111;
        r_rabbitpic[1539] <= 4'b1111;
        r_rabbitpic[1540] <= 4'b1111;
        r_rabbitpic[1541] <= 4'b1111;
        r_rabbitpic[1542] <= 4'b1111;
        r_rabbitpic[1543] <= 4'b1111;
        r_rabbitpic[1544] <= 4'b1111;
        r_rabbitpic[1545] <= 4'b1111;
        r_rabbitpic[1546] <= 4'b1111;
        r_rabbitpic[1547] <= 4'b1111;
        r_rabbitpic[1548] <= 4'b1111;
        r_rabbitpic[1549] <= 4'b1111;
        r_rabbitpic[1550] <= 4'b1111;
        r_rabbitpic[1551] <= 4'b1111;
        r_rabbitpic[1552] <= 4'b1111;
        r_rabbitpic[1553] <= 4'b1111;
        r_rabbitpic[1554] <= 4'b1111;
        r_rabbitpic[1555] <= 4'b1111;
        r_rabbitpic[1556] <= 4'b1111;
        r_rabbitpic[1557] <= 4'b1111;
        r_rabbitpic[1558] <= 4'b0000;
        r_rabbitpic[1559] <= 4'b1111;
        r_rabbitpic[1560] <= 4'b1111;
        r_rabbitpic[1561] <= 4'b1111;
        r_rabbitpic[1562] <= 4'b1111;
        r_rabbitpic[1563] <= 4'b1111;
        r_rabbitpic[1564] <= 4'b1111;
        r_rabbitpic[1565] <= 4'b1111;
        r_rabbitpic[1566] <= 4'b1111;
        r_rabbitpic[1567] <= 4'b1111;
        r_rabbitpic[1568] <= 4'b1111;
        r_rabbitpic[1569] <= 4'b1111;
        r_rabbitpic[1570] <= 4'b1111;
        r_rabbitpic[1571] <= 4'b1111;
        r_rabbitpic[1572] <= 4'b1111;
        r_rabbitpic[1573] <= 4'b1111;
        r_rabbitpic[1574] <= 4'b0000;
        r_rabbitpic[1575] <= 4'b0000;
        r_rabbitpic[1576] <= 4'b1111;
        r_rabbitpic[1577] <= 4'b1111;
        r_rabbitpic[1578] <= 4'b1111;
        r_rabbitpic[1579] <= 4'b1111;
        r_rabbitpic[1580] <= 4'b1111;
        r_rabbitpic[1581] <= 4'b1111;
        r_rabbitpic[1582] <= 4'b1111;
        r_rabbitpic[1583] <= 4'b1111;
        r_rabbitpic[1584] <= 4'b1111;
        r_rabbitpic[1585] <= 4'b1111;
        r_rabbitpic[1586] <= 4'b1111;
        r_rabbitpic[1587] <= 4'b1111;
        r_rabbitpic[1588] <= 4'b1111;
        r_rabbitpic[1589] <= 4'b1111;
        r_rabbitpic[1590] <= 4'b1111;
        r_rabbitpic[1591] <= 4'b1111;
        r_rabbitpic[1592] <= 4'b1111;
        r_rabbitpic[1593] <= 4'b1111;
        r_rabbitpic[1594] <= 4'b1111;
        r_rabbitpic[1595] <= 4'b1111;
        r_rabbitpic[1596] <= 4'b1111;
        r_rabbitpic[1597] <= 4'b1111;
        r_rabbitpic[1598] <= 4'b1111;
        r_rabbitpic[1599] <= 4'b1111;
        r_rabbitpic[1600] <= 4'b1111;
        r_rabbitpic[1601] <= 4'b1111;
        r_rabbitpic[1602] <= 4'b1111;
        r_rabbitpic[1603] <= 4'b1111;
        r_rabbitpic[1604] <= 4'b1111;
        r_rabbitpic[1605] <= 4'b1111;
        r_rabbitpic[1606] <= 4'b1111;
        r_rabbitpic[1607] <= 4'b1111;
        r_rabbitpic[1608] <= 4'b1111;
        r_rabbitpic[1609] <= 4'b1111;
        r_rabbitpic[1610] <= 4'b1111;
        r_rabbitpic[1611] <= 4'b1111;
        r_rabbitpic[1612] <= 4'b1111;
        r_rabbitpic[1613] <= 4'b1111;
        r_rabbitpic[1614] <= 4'b1111;
        r_rabbitpic[1615] <= 4'b1111;
        r_rabbitpic[1616] <= 4'b1111;
        r_rabbitpic[1617] <= 4'b1111;
        r_rabbitpic[1618] <= 4'b1111;
        r_rabbitpic[1619] <= 4'b1111;
        r_rabbitpic[1620] <= 4'b1111;
        r_rabbitpic[1621] <= 4'b1111;
        r_rabbitpic[1622] <= 4'b1111;
        r_rabbitpic[1623] <= 4'b1111;
        r_rabbitpic[1624] <= 4'b1111;
        r_rabbitpic[1625] <= 4'b1111;
        r_rabbitpic[1626] <= 4'b1111;
        r_rabbitpic[1627] <= 4'b1111;
        r_rabbitpic[1628] <= 4'b1111;
        r_rabbitpic[1629] <= 4'b1111;
        r_rabbitpic[1630] <= 4'b1111;
        r_rabbitpic[1631] <= 4'b0000;
        r_rabbitpic[1632] <= 4'b0000;
        r_rabbitpic[1633] <= 4'b1111;
        r_rabbitpic[1634] <= 4'b1111;
        r_rabbitpic[1635] <= 4'b1111;
        r_rabbitpic[1636] <= 4'b1111;
        r_rabbitpic[1637] <= 4'b1111;
        r_rabbitpic[1638] <= 4'b1111;
        r_rabbitpic[1639] <= 4'b1111;
        r_rabbitpic[1640] <= 4'b1111;
        r_rabbitpic[1641] <= 4'b1111;
        r_rabbitpic[1642] <= 4'b1111;
        r_rabbitpic[1643] <= 4'b1111;
        r_rabbitpic[1644] <= 4'b1111;
        r_rabbitpic[1645] <= 4'b1111;
        r_rabbitpic[1646] <= 4'b1111;
        r_rabbitpic[1647] <= 4'b1111;
        r_rabbitpic[1648] <= 4'b1111;
        r_rabbitpic[1649] <= 4'b1111;
        r_rabbitpic[1650] <= 4'b1111;
        r_rabbitpic[1651] <= 4'b1111;
        r_rabbitpic[1652] <= 4'b1111;
        r_rabbitpic[1653] <= 4'b1111;
        r_rabbitpic[1654] <= 4'b1111;
        r_rabbitpic[1655] <= 4'b1111;
        r_rabbitpic[1656] <= 4'b1111;
        r_rabbitpic[1657] <= 4'b1111;
        r_rabbitpic[1658] <= 4'b1111;
        r_rabbitpic[1659] <= 4'b1111;
        r_rabbitpic[1660] <= 4'b1111;
        r_rabbitpic[1661] <= 4'b1111;
        r_rabbitpic[1662] <= 4'b1111;
        r_rabbitpic[1663] <= 4'b1111;
        r_rabbitpic[1664] <= 4'b1111;
        r_rabbitpic[1665] <= 4'b1111;
        r_rabbitpic[1666] <= 4'b1111;
        r_rabbitpic[1667] <= 4'b1111;
        r_rabbitpic[1668] <= 4'b1111;
        r_rabbitpic[1669] <= 4'b1111;
        r_rabbitpic[1670] <= 4'b1111;
        r_rabbitpic[1671] <= 4'b1111;
        r_rabbitpic[1672] <= 4'b1111;
        r_rabbitpic[1673] <= 4'b1111;
        r_rabbitpic[1674] <= 4'b1111;
        r_rabbitpic[1675] <= 4'b1111;
        r_rabbitpic[1676] <= 4'b1111;
        r_rabbitpic[1677] <= 4'b1111;
        r_rabbitpic[1678] <= 4'b1111;
        r_rabbitpic[1679] <= 4'b1111;
        r_rabbitpic[1680] <= 4'b1111;
        r_rabbitpic[1681] <= 4'b1111;
        r_rabbitpic[1682] <= 4'b1111;
        r_rabbitpic[1683] <= 4'b1111;
        r_rabbitpic[1684] <= 4'b1111;
        r_rabbitpic[1685] <= 4'b1111;
        r_rabbitpic[1686] <= 4'b1111;
        r_rabbitpic[1687] <= 4'b0000;
        r_rabbitpic[1688] <= 4'b0000;
        r_rabbitpic[1689] <= 4'b1111;
        r_rabbitpic[1690] <= 4'b1111;
        r_rabbitpic[1691] <= 4'b1111;
        r_rabbitpic[1692] <= 4'b1111;
        r_rabbitpic[1693] <= 4'b1111;
        r_rabbitpic[1694] <= 4'b1111;
        r_rabbitpic[1695] <= 4'b1111;
        r_rabbitpic[1696] <= 4'b1111;
        r_rabbitpic[1697] <= 4'b1111;
        r_rabbitpic[1698] <= 4'b1111;
        r_rabbitpic[1699] <= 4'b1111;
        r_rabbitpic[1700] <= 4'b1111;
        r_rabbitpic[1701] <= 4'b1111;
        r_rabbitpic[1702] <= 4'b1111;
        r_rabbitpic[1703] <= 4'b1111;
        r_rabbitpic[1704] <= 4'b1111;
        r_rabbitpic[1705] <= 4'b1111;
        r_rabbitpic[1706] <= 4'b1111;
        r_rabbitpic[1707] <= 4'b1111;
        r_rabbitpic[1708] <= 4'b1111;
        r_rabbitpic[1709] <= 4'b1111;
        r_rabbitpic[1710] <= 4'b1111;
        r_rabbitpic[1711] <= 4'b1111;
        r_rabbitpic[1712] <= 4'b1111;
        r_rabbitpic[1713] <= 4'b1111;
        r_rabbitpic[1714] <= 4'b1111;
        r_rabbitpic[1715] <= 4'b1111;
        r_rabbitpic[1716] <= 4'b1111;
        r_rabbitpic[1717] <= 4'b1111;
        r_rabbitpic[1718] <= 4'b1111;
        r_rabbitpic[1719] <= 4'b1111;
        r_rabbitpic[1720] <= 4'b1111;
        r_rabbitpic[1721] <= 4'b1111;
        r_rabbitpic[1722] <= 4'b1111;
        r_rabbitpic[1723] <= 4'b1111;
        r_rabbitpic[1724] <= 4'b1111;
        r_rabbitpic[1725] <= 4'b1111;
        r_rabbitpic[1726] <= 4'b1111;
        r_rabbitpic[1727] <= 4'b1111;
        r_rabbitpic[1728] <= 4'b1111;
        r_rabbitpic[1729] <= 4'b1111;
        r_rabbitpic[1730] <= 4'b1111;
        r_rabbitpic[1731] <= 4'b1111;
        r_rabbitpic[1732] <= 4'b1111;
        r_rabbitpic[1733] <= 4'b1111;
        r_rabbitpic[1734] <= 4'b1111;
        r_rabbitpic[1735] <= 4'b1111;
        r_rabbitpic[1736] <= 4'b1111;
        r_rabbitpic[1737] <= 4'b1111;
        r_rabbitpic[1738] <= 4'b1111;
        r_rabbitpic[1739] <= 4'b1111;
        r_rabbitpic[1740] <= 4'b1111;
        r_rabbitpic[1741] <= 4'b1111;
        r_rabbitpic[1742] <= 4'b1111;
        r_rabbitpic[1743] <= 4'b1111;
        r_rabbitpic[1744] <= 4'b0000;
        r_rabbitpic[1745] <= 4'b1111;
        r_rabbitpic[1746] <= 4'b1111;
        r_rabbitpic[1747] <= 4'b1111;
        r_rabbitpic[1748] <= 4'b1111;
        r_rabbitpic[1749] <= 4'b1111;
        r_rabbitpic[1750] <= 4'b1111;
        r_rabbitpic[1751] <= 4'b1111;
        r_rabbitpic[1752] <= 4'b1111;
        r_rabbitpic[1753] <= 4'b1111;
        r_rabbitpic[1754] <= 4'b1111;
        r_rabbitpic[1755] <= 4'b1111;
        r_rabbitpic[1756] <= 4'b1111;
        r_rabbitpic[1757] <= 4'b1111;
        r_rabbitpic[1758] <= 4'b1111;
        r_rabbitpic[1759] <= 4'b1111;
        r_rabbitpic[1760] <= 4'b1111;
        r_rabbitpic[1761] <= 4'b1111;
        r_rabbitpic[1762] <= 4'b1111;
        r_rabbitpic[1763] <= 4'b1111;
        r_rabbitpic[1764] <= 4'b1111;
        r_rabbitpic[1765] <= 4'b1111;
        r_rabbitpic[1766] <= 4'b1111;
        r_rabbitpic[1767] <= 4'b1111;
        r_rabbitpic[1768] <= 4'b1111;
        r_rabbitpic[1769] <= 4'b1111;
        r_rabbitpic[1770] <= 4'b1111;
        r_rabbitpic[1771] <= 4'b1111;
        r_rabbitpic[1772] <= 4'b1111;
        r_rabbitpic[1773] <= 4'b1111;
        r_rabbitpic[1774] <= 4'b1111;
        r_rabbitpic[1775] <= 4'b1111;
        r_rabbitpic[1776] <= 4'b1111;
        r_rabbitpic[1777] <= 4'b1111;
        r_rabbitpic[1778] <= 4'b0000;
        r_rabbitpic[1779] <= 4'b1111;
        r_rabbitpic[1780] <= 4'b1111;
        r_rabbitpic[1781] <= 4'b1111;
        r_rabbitpic[1782] <= 4'b1111;
        r_rabbitpic[1783] <= 4'b1111;
        r_rabbitpic[1784] <= 4'b1111;
        r_rabbitpic[1785] <= 4'b1111;
        r_rabbitpic[1786] <= 4'b1111;
        r_rabbitpic[1787] <= 4'b1111;
        r_rabbitpic[1788] <= 4'b1111;
        r_rabbitpic[1789] <= 4'b1111;
        r_rabbitpic[1790] <= 4'b1111;
        r_rabbitpic[1791] <= 4'b1111;
        r_rabbitpic[1792] <= 4'b1111;
        r_rabbitpic[1793] <= 4'b1111;
        r_rabbitpic[1794] <= 4'b1111;
        r_rabbitpic[1795] <= 4'b1111;
        r_rabbitpic[1796] <= 4'b1111;
        r_rabbitpic[1797] <= 4'b1111;
        r_rabbitpic[1798] <= 4'b1111;
        r_rabbitpic[1799] <= 4'b1111;
        r_rabbitpic[1800] <= 4'b0000;
        r_rabbitpic[1801] <= 4'b1111;
        r_rabbitpic[1802] <= 4'b1111;
        r_rabbitpic[1803] <= 4'b1111;
        r_rabbitpic[1804] <= 4'b1111;
        r_rabbitpic[1805] <= 4'b1111;
        r_rabbitpic[1806] <= 4'b1111;
        r_rabbitpic[1807] <= 4'b1111;
        r_rabbitpic[1808] <= 4'b1111;
        r_rabbitpic[1809] <= 4'b1111;
        r_rabbitpic[1810] <= 4'b1111;
        r_rabbitpic[1811] <= 4'b1111;
        r_rabbitpic[1812] <= 4'b1111;
        r_rabbitpic[1813] <= 4'b1111;
        r_rabbitpic[1814] <= 4'b1111;
        r_rabbitpic[1815] <= 4'b1111;
        r_rabbitpic[1816] <= 4'b1111;
        r_rabbitpic[1817] <= 4'b1111;
        r_rabbitpic[1818] <= 4'b1111;
        r_rabbitpic[1819] <= 4'b1111;
        r_rabbitpic[1820] <= 4'b1111;
        r_rabbitpic[1821] <= 4'b1111;
        r_rabbitpic[1822] <= 4'b1111;
        r_rabbitpic[1823] <= 4'b1111;
        r_rabbitpic[1824] <= 4'b1111;
        r_rabbitpic[1825] <= 4'b1111;
        r_rabbitpic[1826] <= 4'b1111;
        r_rabbitpic[1827] <= 4'b1111;
        r_rabbitpic[1828] <= 4'b1111;
        r_rabbitpic[1829] <= 4'b1111;
        r_rabbitpic[1830] <= 4'b1111;
        r_rabbitpic[1831] <= 4'b1111;
        r_rabbitpic[1832] <= 4'b1111;
        r_rabbitpic[1833] <= 4'b0000;
        r_rabbitpic[1834] <= 4'b1111;
        r_rabbitpic[1835] <= 4'b0000;
        r_rabbitpic[1836] <= 4'b1111;
        r_rabbitpic[1837] <= 4'b1111;
        r_rabbitpic[1838] <= 4'b1111;
        r_rabbitpic[1839] <= 4'b1111;
        r_rabbitpic[1840] <= 4'b1111;
        r_rabbitpic[1841] <= 4'b1111;
        r_rabbitpic[1842] <= 4'b1111;
        r_rabbitpic[1843] <= 4'b1111;
        r_rabbitpic[1844] <= 4'b1111;
        r_rabbitpic[1845] <= 4'b1111;
        r_rabbitpic[1846] <= 4'b1111;
        r_rabbitpic[1847] <= 4'b1111;
        r_rabbitpic[1848] <= 4'b1111;
        r_rabbitpic[1849] <= 4'b1111;
        r_rabbitpic[1850] <= 4'b1111;
        r_rabbitpic[1851] <= 4'b1111;
        r_rabbitpic[1852] <= 4'b1111;
        r_rabbitpic[1853] <= 4'b1111;
        r_rabbitpic[1854] <= 4'b1111;
        r_rabbitpic[1855] <= 4'b0000;
        r_rabbitpic[1856] <= 4'b1111;
        r_rabbitpic[1857] <= 4'b1111;
        r_rabbitpic[1858] <= 4'b1111;
        r_rabbitpic[1859] <= 4'b1111;
        r_rabbitpic[1860] <= 4'b1111;
        r_rabbitpic[1861] <= 4'b1111;
        r_rabbitpic[1862] <= 4'b1111;
        r_rabbitpic[1863] <= 4'b1111;
        r_rabbitpic[1864] <= 4'b1111;
        r_rabbitpic[1865] <= 4'b1111;
        r_rabbitpic[1866] <= 4'b1111;
        r_rabbitpic[1867] <= 4'b1111;
        r_rabbitpic[1868] <= 4'b1111;
        r_rabbitpic[1869] <= 4'b1111;
        r_rabbitpic[1870] <= 4'b1111;
        r_rabbitpic[1871] <= 4'b1111;
        r_rabbitpic[1872] <= 4'b1111;
        r_rabbitpic[1873] <= 4'b1111;
        r_rabbitpic[1874] <= 4'b1111;
        r_rabbitpic[1875] <= 4'b1111;
        r_rabbitpic[1876] <= 4'b1111;
        r_rabbitpic[1877] <= 4'b1111;
        r_rabbitpic[1878] <= 4'b1111;
        r_rabbitpic[1879] <= 4'b1111;
        r_rabbitpic[1880] <= 4'b1111;
        r_rabbitpic[1881] <= 4'b1111;
        r_rabbitpic[1882] <= 4'b1111;
        r_rabbitpic[1883] <= 4'b1111;
        r_rabbitpic[1884] <= 4'b1111;
        r_rabbitpic[1885] <= 4'b1111;
        r_rabbitpic[1886] <= 4'b1111;
        r_rabbitpic[1887] <= 4'b1111;
        r_rabbitpic[1888] <= 4'b0000;
        r_rabbitpic[1889] <= 4'b0000;
        r_rabbitpic[1890] <= 4'b0000;
        r_rabbitpic[1891] <= 4'b1111;
        r_rabbitpic[1892] <= 4'b1111;
        r_rabbitpic[1893] <= 4'b1111;
        r_rabbitpic[1894] <= 4'b1111;
        r_rabbitpic[1895] <= 4'b1111;
        r_rabbitpic[1896] <= 4'b1111;
        r_rabbitpic[1897] <= 4'b1111;
        r_rabbitpic[1898] <= 4'b1111;
        r_rabbitpic[1899] <= 4'b1111;
        r_rabbitpic[1900] <= 4'b1111;
        r_rabbitpic[1901] <= 4'b1111;
        r_rabbitpic[1902] <= 4'b1111;
        r_rabbitpic[1903] <= 4'b1111;
        r_rabbitpic[1904] <= 4'b1111;
        r_rabbitpic[1905] <= 4'b0000;
        r_rabbitpic[1906] <= 4'b0000;
        r_rabbitpic[1907] <= 4'b1111;
        r_rabbitpic[1908] <= 4'b1111;
        r_rabbitpic[1909] <= 4'b1111;
        r_rabbitpic[1910] <= 4'b1111;
        r_rabbitpic[1911] <= 4'b0000;
        r_rabbitpic[1912] <= 4'b1111;
        r_rabbitpic[1913] <= 4'b1111;
        r_rabbitpic[1914] <= 4'b1111;
        r_rabbitpic[1915] <= 4'b1111;
        r_rabbitpic[1916] <= 4'b1111;
        r_rabbitpic[1917] <= 4'b1111;
        r_rabbitpic[1918] <= 4'b1111;
        r_rabbitpic[1919] <= 4'b1111;
        r_rabbitpic[1920] <= 4'b1111;
        r_rabbitpic[1921] <= 4'b1111;
        r_rabbitpic[1922] <= 4'b1111;
        r_rabbitpic[1923] <= 4'b1111;
        r_rabbitpic[1924] <= 4'b1111;
        r_rabbitpic[1925] <= 4'b1111;
        r_rabbitpic[1926] <= 4'b1111;
        r_rabbitpic[1927] <= 4'b1111;
        r_rabbitpic[1928] <= 4'b1111;
        r_rabbitpic[1929] <= 4'b1111;
        r_rabbitpic[1930] <= 4'b1111;
        r_rabbitpic[1931] <= 4'b1111;
        r_rabbitpic[1932] <= 4'b1111;
        r_rabbitpic[1933] <= 4'b1111;
        r_rabbitpic[1934] <= 4'b1111;
        r_rabbitpic[1935] <= 4'b1111;
        r_rabbitpic[1936] <= 4'b1111;
        r_rabbitpic[1937] <= 4'b1111;
        r_rabbitpic[1938] <= 4'b1111;
        r_rabbitpic[1939] <= 4'b1111;
        r_rabbitpic[1940] <= 4'b0000;
        r_rabbitpic[1941] <= 4'b0000;
        r_rabbitpic[1942] <= 4'b0000;
        r_rabbitpic[1943] <= 4'b1111;
        r_rabbitpic[1944] <= 4'b0000;
        r_rabbitpic[1945] <= 4'b0000;
        r_rabbitpic[1946] <= 4'b1111;
        r_rabbitpic[1947] <= 4'b1111;
        r_rabbitpic[1948] <= 4'b1111;
        r_rabbitpic[1949] <= 4'b1111;
        r_rabbitpic[1950] <= 4'b1111;
        r_rabbitpic[1951] <= 4'b1111;
        r_rabbitpic[1952] <= 4'b1111;
        r_rabbitpic[1953] <= 4'b1111;
        r_rabbitpic[1954] <= 4'b1111;
        r_rabbitpic[1955] <= 4'b1111;
        r_rabbitpic[1956] <= 4'b1111;
        r_rabbitpic[1957] <= 4'b1111;
        r_rabbitpic[1958] <= 4'b1111;
        r_rabbitpic[1959] <= 4'b0000;
        r_rabbitpic[1960] <= 4'b1111;
        r_rabbitpic[1961] <= 4'b1111;
        r_rabbitpic[1962] <= 4'b1111;
        r_rabbitpic[1963] <= 4'b1111;
        r_rabbitpic[1964] <= 4'b1111;
        r_rabbitpic[1965] <= 4'b1111;
        r_rabbitpic[1966] <= 4'b0000;
        r_rabbitpic[1967] <= 4'b1111;
        r_rabbitpic[1968] <= 4'b1111;
        r_rabbitpic[1969] <= 4'b1111;
        r_rabbitpic[1970] <= 4'b1111;
        r_rabbitpic[1971] <= 4'b1111;
        r_rabbitpic[1972] <= 4'b1111;
        r_rabbitpic[1973] <= 4'b1111;
        r_rabbitpic[1974] <= 4'b1111;
        r_rabbitpic[1975] <= 4'b1111;
        r_rabbitpic[1976] <= 4'b1111;
        r_rabbitpic[1977] <= 4'b1111;
        r_rabbitpic[1978] <= 4'b1111;
        r_rabbitpic[1979] <= 4'b1111;
        r_rabbitpic[1980] <= 4'b1111;
        r_rabbitpic[1981] <= 4'b1111;
        r_rabbitpic[1982] <= 4'b1111;
        r_rabbitpic[1983] <= 4'b1111;
        r_rabbitpic[1984] <= 4'b1111;
        r_rabbitpic[1985] <= 4'b1111;
        r_rabbitpic[1986] <= 4'b1111;
        r_rabbitpic[1987] <= 4'b1111;
        r_rabbitpic[1988] <= 4'b1111;
        r_rabbitpic[1989] <= 4'b1111;
        r_rabbitpic[1990] <= 4'b1111;
        r_rabbitpic[1991] <= 4'b1111;
        r_rabbitpic[1992] <= 4'b1111;
        r_rabbitpic[1993] <= 4'b1111;
        r_rabbitpic[1994] <= 4'b0000;
        r_rabbitpic[1995] <= 4'b1111;
        r_rabbitpic[1996] <= 4'b1111;
        r_rabbitpic[1997] <= 4'b1111;
        r_rabbitpic[1998] <= 4'b0000;
        r_rabbitpic[1999] <= 4'b0000;
        r_rabbitpic[2000] <= 4'b0000;
        r_rabbitpic[2001] <= 4'b0000;
        r_rabbitpic[2002] <= 4'b1111;
        r_rabbitpic[2003] <= 4'b1111;
        r_rabbitpic[2004] <= 4'b1111;
        r_rabbitpic[2005] <= 4'b1111;
        r_rabbitpic[2006] <= 4'b1111;
        r_rabbitpic[2007] <= 4'b0000;
        r_rabbitpic[2008] <= 4'b1111;
        r_rabbitpic[2009] <= 4'b1111;
        r_rabbitpic[2010] <= 4'b1111;
        r_rabbitpic[2011] <= 4'b1111;
        r_rabbitpic[2012] <= 4'b1111;
        r_rabbitpic[2013] <= 4'b0000;
        r_rabbitpic[2014] <= 4'b1111;
        r_rabbitpic[2015] <= 4'b1111;
        r_rabbitpic[2016] <= 4'b1111;
        r_rabbitpic[2017] <= 4'b1111;
        r_rabbitpic[2018] <= 4'b1111;
        r_rabbitpic[2019] <= 4'b1111;
        r_rabbitpic[2020] <= 4'b1111;
        r_rabbitpic[2021] <= 4'b1111;
        r_rabbitpic[2022] <= 4'b0000;
        r_rabbitpic[2023] <= 4'b1111;
        r_rabbitpic[2024] <= 4'b1111;
        r_rabbitpic[2025] <= 4'b1111;
        r_rabbitpic[2026] <= 4'b1111;
        r_rabbitpic[2027] <= 4'b1111;
        r_rabbitpic[2028] <= 4'b1111;
        r_rabbitpic[2029] <= 4'b1111;
        r_rabbitpic[2030] <= 4'b1111;
        r_rabbitpic[2031] <= 4'b1111;
        r_rabbitpic[2032] <= 4'b1111;
        r_rabbitpic[2033] <= 4'b1111;
        r_rabbitpic[2034] <= 4'b1111;
        r_rabbitpic[2035] <= 4'b1111;
        r_rabbitpic[2036] <= 4'b1111;
        r_rabbitpic[2037] <= 4'b1111;
        r_rabbitpic[2038] <= 4'b1111;
        r_rabbitpic[2039] <= 4'b1111;
        r_rabbitpic[2040] <= 4'b1111;
        r_rabbitpic[2041] <= 4'b1111;
        r_rabbitpic[2042] <= 4'b1111;
        r_rabbitpic[2043] <= 4'b1111;
        r_rabbitpic[2044] <= 4'b1111;
        r_rabbitpic[2045] <= 4'b1111;
        r_rabbitpic[2046] <= 4'b1111;
        r_rabbitpic[2047] <= 4'b1111;
        r_rabbitpic[2048] <= 4'b1111;
        r_rabbitpic[2049] <= 4'b0000;
        r_rabbitpic[2050] <= 4'b1111;
        r_rabbitpic[2051] <= 4'b1111;
        r_rabbitpic[2052] <= 4'b1111;
        r_rabbitpic[2053] <= 4'b1111;
        r_rabbitpic[2054] <= 4'b1111;
        r_rabbitpic[2055] <= 4'b1111;
        r_rabbitpic[2056] <= 4'b0000;
        r_rabbitpic[2057] <= 4'b1111;
        r_rabbitpic[2058] <= 4'b1111;
        r_rabbitpic[2059] <= 4'b1111;
        r_rabbitpic[2060] <= 4'b1111;
        r_rabbitpic[2061] <= 4'b0000;
        r_rabbitpic[2062] <= 4'b1111;
        r_rabbitpic[2063] <= 4'b1111;
        r_rabbitpic[2064] <= 4'b0000;
        r_rabbitpic[2065] <= 4'b0000;
        r_rabbitpic[2066] <= 4'b1111;
        r_rabbitpic[2067] <= 4'b1111;
        r_rabbitpic[2068] <= 4'b1111;
        r_rabbitpic[2069] <= 4'b1111;
        r_rabbitpic[2070] <= 4'b1111;
        r_rabbitpic[2071] <= 4'b1111;
        r_rabbitpic[2072] <= 4'b1111;
        r_rabbitpic[2073] <= 4'b1111;
        r_rabbitpic[2074] <= 4'b1111;
        r_rabbitpic[2075] <= 4'b1111;
        r_rabbitpic[2076] <= 4'b1111;
        r_rabbitpic[2077] <= 4'b0000;
        r_rabbitpic[2078] <= 4'b1111;
        r_rabbitpic[2079] <= 4'b1111;
        r_rabbitpic[2080] <= 4'b1111;
        r_rabbitpic[2081] <= 4'b1111;
        r_rabbitpic[2082] <= 4'b1111;
        r_rabbitpic[2083] <= 4'b1111;
        r_rabbitpic[2084] <= 4'b1111;
        r_rabbitpic[2085] <= 4'b1111;
        r_rabbitpic[2086] <= 4'b1111;
        r_rabbitpic[2087] <= 4'b1111;
        r_rabbitpic[2088] <= 4'b1111;
        r_rabbitpic[2089] <= 4'b1111;
        r_rabbitpic[2090] <= 4'b1111;
        r_rabbitpic[2091] <= 4'b1111;
        r_rabbitpic[2092] <= 4'b1111;
        r_rabbitpic[2093] <= 4'b1111;
        r_rabbitpic[2094] <= 4'b1111;
        r_rabbitpic[2095] <= 4'b1111;
        r_rabbitpic[2096] <= 4'b1111;
        r_rabbitpic[2097] <= 4'b1111;
        r_rabbitpic[2098] <= 4'b1111;
        r_rabbitpic[2099] <= 4'b1111;
        r_rabbitpic[2100] <= 4'b1111;
        r_rabbitpic[2101] <= 4'b1111;
        r_rabbitpic[2102] <= 4'b1111;
        r_rabbitpic[2103] <= 4'b0000;
        r_rabbitpic[2104] <= 4'b1111;
        r_rabbitpic[2105] <= 4'b0000;
        r_rabbitpic[2106] <= 4'b1111;
        r_rabbitpic[2107] <= 4'b0000;
        r_rabbitpic[2108] <= 4'b0000;
        r_rabbitpic[2109] <= 4'b1111;
        r_rabbitpic[2110] <= 4'b1111;
        r_rabbitpic[2111] <= 4'b1111;
        r_rabbitpic[2112] <= 4'b0000;
        r_rabbitpic[2113] <= 4'b1111;
        r_rabbitpic[2114] <= 4'b1111;
        r_rabbitpic[2115] <= 4'b1111;
        r_rabbitpic[2116] <= 4'b0000;
        r_rabbitpic[2117] <= 4'b1111;
        r_rabbitpic[2118] <= 4'b1111;
        r_rabbitpic[2119] <= 4'b1111;
        r_rabbitpic[2120] <= 4'b1111;
        r_rabbitpic[2121] <= 4'b1111;
        r_rabbitpic[2122] <= 4'b0000;
        r_rabbitpic[2123] <= 4'b1111;
        r_rabbitpic[2124] <= 4'b1111;
        r_rabbitpic[2125] <= 4'b1111;
        r_rabbitpic[2126] <= 4'b1111;
        r_rabbitpic[2127] <= 4'b1111;
        r_rabbitpic[2128] <= 4'b1111;
        r_rabbitpic[2129] <= 4'b1111;
        r_rabbitpic[2130] <= 4'b1111;
        r_rabbitpic[2131] <= 4'b1111;
        r_rabbitpic[2132] <= 4'b1111;
        r_rabbitpic[2133] <= 4'b1111;
        r_rabbitpic[2134] <= 4'b1111;
        r_rabbitpic[2135] <= 4'b1111;
        r_rabbitpic[2136] <= 4'b1111;
        r_rabbitpic[2137] <= 4'b1111;
        r_rabbitpic[2138] <= 4'b1111;
        r_rabbitpic[2139] <= 4'b1111;
        r_rabbitpic[2140] <= 4'b1111;
        r_rabbitpic[2141] <= 4'b1111;
        r_rabbitpic[2142] <= 4'b1111;
        r_rabbitpic[2143] <= 4'b1111;
        r_rabbitpic[2144] <= 4'b1111;
        r_rabbitpic[2145] <= 4'b1111;
        r_rabbitpic[2146] <= 4'b1111;
        r_rabbitpic[2147] <= 4'b1111;
        r_rabbitpic[2148] <= 4'b1111;
        r_rabbitpic[2149] <= 4'b1111;
        r_rabbitpic[2150] <= 4'b1111;
        r_rabbitpic[2151] <= 4'b1111;
        r_rabbitpic[2152] <= 4'b1111;
        r_rabbitpic[2153] <= 4'b1111;
        r_rabbitpic[2154] <= 4'b1111;
        r_rabbitpic[2155] <= 4'b1111;
        r_rabbitpic[2156] <= 4'b1111;
        r_rabbitpic[2157] <= 4'b1111;
        r_rabbitpic[2158] <= 4'b0000;
        r_rabbitpic[2159] <= 4'b1111;
        r_rabbitpic[2160] <= 4'b0000;
        r_rabbitpic[2161] <= 4'b0000;
        r_rabbitpic[2162] <= 4'b0000;
        r_rabbitpic[2163] <= 4'b1111;
        r_rabbitpic[2164] <= 4'b0000;
        r_rabbitpic[2165] <= 4'b0000;
        r_rabbitpic[2166] <= 4'b0000;
        r_rabbitpic[2167] <= 4'b0000;
        r_rabbitpic[2168] <= 4'b1111;
        r_rabbitpic[2169] <= 4'b1111;
        r_rabbitpic[2170] <= 4'b0000;
        r_rabbitpic[2171] <= 4'b0000;
        r_rabbitpic[2172] <= 4'b1111;
        r_rabbitpic[2173] <= 4'b1111;
        r_rabbitpic[2174] <= 4'b1111;
        r_rabbitpic[2175] <= 4'b1111;
        r_rabbitpic[2176] <= 4'b1111;
        r_rabbitpic[2177] <= 4'b0000;
        r_rabbitpic[2178] <= 4'b1111;
        r_rabbitpic[2179] <= 4'b1111;
        r_rabbitpic[2180] <= 4'b1111;
        r_rabbitpic[2181] <= 4'b1111;
        r_rabbitpic[2182] <= 4'b1111;
        r_rabbitpic[2183] <= 4'b1111;
        r_rabbitpic[2184] <= 4'b1111;
        r_rabbitpic[2185] <= 4'b1111;
        r_rabbitpic[2186] <= 4'b1111;
        r_rabbitpic[2187] <= 4'b1111;
        r_rabbitpic[2188] <= 4'b0000;
        r_rabbitpic[2189] <= 4'b0000;
        r_rabbitpic[2190] <= 4'b1111;
        r_rabbitpic[2191] <= 4'b1111;
        r_rabbitpic[2192] <= 4'b1111;
        r_rabbitpic[2193] <= 4'b1111;
        r_rabbitpic[2194] <= 4'b1111;
        r_rabbitpic[2195] <= 4'b1111;
        r_rabbitpic[2196] <= 4'b1111;
        r_rabbitpic[2197] <= 4'b1111;
        r_rabbitpic[2198] <= 4'b1111;
        r_rabbitpic[2199] <= 4'b1111;
        r_rabbitpic[2200] <= 4'b1111;
        r_rabbitpic[2201] <= 4'b1111;
        r_rabbitpic[2202] <= 4'b1111;
        r_rabbitpic[2203] <= 4'b1111;
        r_rabbitpic[2204] <= 4'b1111;
        r_rabbitpic[2205] <= 4'b1111;
        r_rabbitpic[2206] <= 4'b1111;
        r_rabbitpic[2207] <= 4'b1111;
        r_rabbitpic[2208] <= 4'b1111;
        r_rabbitpic[2209] <= 4'b1111;
        r_rabbitpic[2210] <= 4'b1111;
        r_rabbitpic[2211] <= 4'b1111;
        r_rabbitpic[2212] <= 4'b1111;
        r_rabbitpic[2213] <= 4'b1111;
        r_rabbitpic[2214] <= 4'b0000;
        r_rabbitpic[2215] <= 4'b0000;
        r_rabbitpic[2216] <= 4'b0000;
        r_rabbitpic[2217] <= 4'b1111;
        r_rabbitpic[2218] <= 4'b1111;
        r_rabbitpic[2219] <= 4'b1111;
        r_rabbitpic[2220] <= 4'b1111;
        r_rabbitpic[2221] <= 4'b0000;
        r_rabbitpic[2222] <= 4'b1111;
        r_rabbitpic[2223] <= 4'b1111;
        r_rabbitpic[2224] <= 4'b0000;
        r_rabbitpic[2225] <= 4'b1111;
        r_rabbitpic[2226] <= 4'b1111;
        r_rabbitpic[2227] <= 4'b0000;
        r_rabbitpic[2228] <= 4'b1111;
        r_rabbitpic[2229] <= 4'b1111;
        r_rabbitpic[2230] <= 4'b1111;
        r_rabbitpic[2231] <= 4'b1111;
        r_rabbitpic[2232] <= 4'b1111;
        r_rabbitpic[2233] <= 4'b0000;
        r_rabbitpic[2234] <= 4'b1111;
        r_rabbitpic[2235] <= 4'b1111;
        r_rabbitpic[2236] <= 4'b1111;
        r_rabbitpic[2237] <= 4'b1111;
        r_rabbitpic[2238] <= 4'b1111;
        r_rabbitpic[2239] <= 4'b1111;
        r_rabbitpic[2240] <= 4'b1111;
        r_rabbitpic[2241] <= 4'b1111;
        r_rabbitpic[2242] <= 4'b1111;
        r_rabbitpic[2243] <= 4'b0000;
        r_rabbitpic[2244] <= 4'b1111;
        r_rabbitpic[2245] <= 4'b0000;
        r_rabbitpic[2246] <= 4'b1111;
        r_rabbitpic[2247] <= 4'b1111;
        r_rabbitpic[2248] <= 4'b1111;
        r_rabbitpic[2249] <= 4'b1111;
        r_rabbitpic[2250] <= 4'b1111;
        r_rabbitpic[2251] <= 4'b1111;
        r_rabbitpic[2252] <= 4'b1111;
        r_rabbitpic[2253] <= 4'b1111;
        r_rabbitpic[2254] <= 4'b1111;
        r_rabbitpic[2255] <= 4'b1111;
        r_rabbitpic[2256] <= 4'b1111;
        r_rabbitpic[2257] <= 4'b1111;
        r_rabbitpic[2258] <= 4'b1111;
        r_rabbitpic[2259] <= 4'b1111;
        r_rabbitpic[2260] <= 4'b1111;
        r_rabbitpic[2261] <= 4'b1111;
        r_rabbitpic[2262] <= 4'b1111;
        r_rabbitpic[2263] <= 4'b1111;
        r_rabbitpic[2264] <= 4'b1111;
        r_rabbitpic[2265] <= 4'b1111;
        r_rabbitpic[2266] <= 4'b1111;
        r_rabbitpic[2267] <= 4'b1111;
        r_rabbitpic[2268] <= 4'b1111;
        r_rabbitpic[2269] <= 4'b1111;
        r_rabbitpic[2270] <= 4'b1111;
        r_rabbitpic[2271] <= 4'b1111;
        r_rabbitpic[2272] <= 4'b1111;
        r_rabbitpic[2273] <= 4'b1111;
        r_rabbitpic[2274] <= 4'b1111;
        r_rabbitpic[2275] <= 4'b1111;
        r_rabbitpic[2276] <= 4'b0000;
        r_rabbitpic[2277] <= 4'b1111;
        r_rabbitpic[2278] <= 4'b1111;
        r_rabbitpic[2279] <= 4'b0000;
        r_rabbitpic[2280] <= 4'b1111;
        r_rabbitpic[2281] <= 4'b1111;
        r_rabbitpic[2282] <= 4'b0000;
        r_rabbitpic[2283] <= 4'b1111;
        r_rabbitpic[2284] <= 4'b1111;
        r_rabbitpic[2285] <= 4'b1111;
        r_rabbitpic[2286] <= 4'b1111;
        r_rabbitpic[2287] <= 4'b1111;
        r_rabbitpic[2288] <= 4'b0000;
        r_rabbitpic[2289] <= 4'b1111;
        r_rabbitpic[2290] <= 4'b1111;
        r_rabbitpic[2291] <= 4'b1111;
        r_rabbitpic[2292] <= 4'b1111;
        r_rabbitpic[2293] <= 4'b1111;
        r_rabbitpic[2294] <= 4'b1111;
        r_rabbitpic[2295] <= 4'b1111;
        r_rabbitpic[2296] <= 4'b1111;
        r_rabbitpic[2297] <= 4'b1111;
        r_rabbitpic[2298] <= 4'b0000;
        r_rabbitpic[2299] <= 4'b1111;
        r_rabbitpic[2300] <= 4'b0000;
        r_rabbitpic[2301] <= 4'b1111;
        r_rabbitpic[2302] <= 4'b1111;
        r_rabbitpic[2303] <= 4'b1111;
        r_rabbitpic[2304] <= 4'b1111;
        r_rabbitpic[2305] <= 4'b1111;
        r_rabbitpic[2306] <= 4'b1111;
        r_rabbitpic[2307] <= 4'b1111;
        r_rabbitpic[2308] <= 4'b1111;
        r_rabbitpic[2309] <= 4'b1111;
        r_rabbitpic[2310] <= 4'b1111;
        r_rabbitpic[2311] <= 4'b1111;
        r_rabbitpic[2312] <= 4'b1111;
        r_rabbitpic[2313] <= 4'b1111;
        r_rabbitpic[2314] <= 4'b1111;
        r_rabbitpic[2315] <= 4'b1111;
        r_rabbitpic[2316] <= 4'b1111;
        r_rabbitpic[2317] <= 4'b1111;
        r_rabbitpic[2318] <= 4'b1111;
        r_rabbitpic[2319] <= 4'b1111;
        r_rabbitpic[2320] <= 4'b1111;
        r_rabbitpic[2321] <= 4'b1111;
        r_rabbitpic[2322] <= 4'b1111;
        r_rabbitpic[2323] <= 4'b1111;
        r_rabbitpic[2324] <= 4'b1111;
        r_rabbitpic[2325] <= 4'b1111;
        r_rabbitpic[2326] <= 4'b1111;
        r_rabbitpic[2327] <= 4'b1111;
        r_rabbitpic[2328] <= 4'b1111;
        r_rabbitpic[2329] <= 4'b1111;
        r_rabbitpic[2330] <= 4'b1111;
        r_rabbitpic[2331] <= 4'b0000;
        r_rabbitpic[2332] <= 4'b1111;
        r_rabbitpic[2333] <= 4'b0000;
        r_rabbitpic[2334] <= 4'b1111;
        r_rabbitpic[2335] <= 4'b1111;
        r_rabbitpic[2336] <= 4'b1111;
        r_rabbitpic[2337] <= 4'b1111;
        r_rabbitpic[2338] <= 4'b0000;
        r_rabbitpic[2339] <= 4'b1111;
        r_rabbitpic[2340] <= 4'b1111;
        r_rabbitpic[2341] <= 4'b1111;
        r_rabbitpic[2342] <= 4'b1111;
        r_rabbitpic[2343] <= 4'b1111;
        r_rabbitpic[2344] <= 4'b0000;
        r_rabbitpic[2345] <= 4'b1111;
        r_rabbitpic[2346] <= 4'b1111;
        r_rabbitpic[2347] <= 4'b1111;
        r_rabbitpic[2348] <= 4'b1111;
        r_rabbitpic[2349] <= 4'b1111;
        r_rabbitpic[2350] <= 4'b1111;
        r_rabbitpic[2351] <= 4'b1111;
        r_rabbitpic[2352] <= 4'b1111;
        r_rabbitpic[2353] <= 4'b0000;
        r_rabbitpic[2354] <= 4'b1111;
        r_rabbitpic[2355] <= 4'b0000;
        r_rabbitpic[2356] <= 4'b1111;
        r_rabbitpic[2357] <= 4'b1111;
        r_rabbitpic[2358] <= 4'b1111;
        r_rabbitpic[2359] <= 4'b1111;
        r_rabbitpic[2360] <= 4'b1111;
        r_rabbitpic[2361] <= 4'b1111;
        r_rabbitpic[2362] <= 4'b1111;
        r_rabbitpic[2363] <= 4'b1111;
        r_rabbitpic[2364] <= 4'b1111;
        r_rabbitpic[2365] <= 4'b1111;
        r_rabbitpic[2366] <= 4'b1111;
        r_rabbitpic[2367] <= 4'b1111;
        r_rabbitpic[2368] <= 4'b1111;
        r_rabbitpic[2369] <= 4'b1111;
        r_rabbitpic[2370] <= 4'b1111;
        r_rabbitpic[2371] <= 4'b1111;
        r_rabbitpic[2372] <= 4'b1111;
        r_rabbitpic[2373] <= 4'b1111;
        r_rabbitpic[2374] <= 4'b1111;
        r_rabbitpic[2375] <= 4'b1111;
        r_rabbitpic[2376] <= 4'b1111;
        r_rabbitpic[2377] <= 4'b1111;
        r_rabbitpic[2378] <= 4'b1111;
        r_rabbitpic[2379] <= 4'b1111;
        r_rabbitpic[2380] <= 4'b1111;
        r_rabbitpic[2381] <= 4'b1111;
        r_rabbitpic[2382] <= 4'b1111;
        r_rabbitpic[2383] <= 4'b1111;
        r_rabbitpic[2384] <= 4'b1111;
        r_rabbitpic[2385] <= 4'b0000;
        r_rabbitpic[2386] <= 4'b1111;
        r_rabbitpic[2387] <= 4'b1111;
        r_rabbitpic[2388] <= 4'b0000;
        r_rabbitpic[2389] <= 4'b1111;
        r_rabbitpic[2390] <= 4'b1111;
        r_rabbitpic[2391] <= 4'b1111;
        r_rabbitpic[2392] <= 4'b1111;
        r_rabbitpic[2393] <= 4'b0000;
        r_rabbitpic[2394] <= 4'b0000;
        r_rabbitpic[2395] <= 4'b1111;
        r_rabbitpic[2396] <= 4'b1111;
        r_rabbitpic[2397] <= 4'b1111;
        r_rabbitpic[2398] <= 4'b1111;
        r_rabbitpic[2399] <= 4'b1111;
        r_rabbitpic[2400] <= 4'b0000;
        r_rabbitpic[2401] <= 4'b1111;
        r_rabbitpic[2402] <= 4'b1111;
        r_rabbitpic[2403] <= 4'b1111;
        r_rabbitpic[2404] <= 4'b1111;
        r_rabbitpic[2405] <= 4'b1111;
        r_rabbitpic[2406] <= 4'b1111;
        r_rabbitpic[2407] <= 4'b0000;
        r_rabbitpic[2408] <= 4'b1111;
        r_rabbitpic[2409] <= 4'b1111;
        r_rabbitpic[2410] <= 4'b0000;
        r_rabbitpic[2411] <= 4'b1111;
        r_rabbitpic[2412] <= 4'b1111;
        r_rabbitpic[2413] <= 4'b1111;
        r_rabbitpic[2414] <= 4'b1111;
        r_rabbitpic[2415] <= 4'b1111;
        r_rabbitpic[2416] <= 4'b1111;
        r_rabbitpic[2417] <= 4'b1111;
        r_rabbitpic[2418] <= 4'b1111;
        r_rabbitpic[2419] <= 4'b1111;
        r_rabbitpic[2420] <= 4'b1111;
        r_rabbitpic[2421] <= 4'b1111;
        r_rabbitpic[2422] <= 4'b1111;
        r_rabbitpic[2423] <= 4'b1111;
        r_rabbitpic[2424] <= 4'b1111;
        r_rabbitpic[2425] <= 4'b1111;
        r_rabbitpic[2426] <= 4'b1111;
        r_rabbitpic[2427] <= 4'b1111;
        r_rabbitpic[2428] <= 4'b1111;
        r_rabbitpic[2429] <= 4'b1111;
        r_rabbitpic[2430] <= 4'b1111;
        r_rabbitpic[2431] <= 4'b1111;
        r_rabbitpic[2432] <= 4'b1111;
        r_rabbitpic[2433] <= 4'b1111;
        r_rabbitpic[2434] <= 4'b1111;
        r_rabbitpic[2435] <= 4'b1111;
        r_rabbitpic[2436] <= 4'b1111;
        r_rabbitpic[2437] <= 4'b1111;
        r_rabbitpic[2438] <= 4'b1111;
        r_rabbitpic[2439] <= 4'b1111;
        r_rabbitpic[2440] <= 4'b0000;
        r_rabbitpic[2441] <= 4'b1111;
        r_rabbitpic[2442] <= 4'b1111;
        r_rabbitpic[2443] <= 4'b0000;
        r_rabbitpic[2444] <= 4'b1111;
        r_rabbitpic[2445] <= 4'b1111;
        r_rabbitpic[2446] <= 4'b1111;
        r_rabbitpic[2447] <= 4'b1111;
        r_rabbitpic[2448] <= 4'b1111;
        r_rabbitpic[2449] <= 4'b0000;
        r_rabbitpic[2450] <= 4'b0000;
        r_rabbitpic[2451] <= 4'b1111;
        r_rabbitpic[2452] <= 4'b1111;
        r_rabbitpic[2453] <= 4'b1111;
        r_rabbitpic[2454] <= 4'b1111;
        r_rabbitpic[2455] <= 4'b1111;
        r_rabbitpic[2456] <= 4'b0000;
        r_rabbitpic[2457] <= 4'b1111;
        r_rabbitpic[2458] <= 4'b1111;
        r_rabbitpic[2459] <= 4'b1111;
        r_rabbitpic[2460] <= 4'b1111;
        r_rabbitpic[2461] <= 4'b1111;
        r_rabbitpic[2462] <= 4'b0000;
        r_rabbitpic[2463] <= 4'b1111;
        r_rabbitpic[2464] <= 4'b1111;
        r_rabbitpic[2465] <= 4'b0000;
        r_rabbitpic[2466] <= 4'b1111;
        r_rabbitpic[2467] <= 4'b1111;
        r_rabbitpic[2468] <= 4'b1111;
        r_rabbitpic[2469] <= 4'b1111;
        r_rabbitpic[2470] <= 4'b1111;
        r_rabbitpic[2471] <= 4'b1111;
        r_rabbitpic[2472] <= 4'b1111;
        r_rabbitpic[2473] <= 4'b1111;
        r_rabbitpic[2474] <= 4'b1111;
        r_rabbitpic[2475] <= 4'b1111;
        r_rabbitpic[2476] <= 4'b1111;
        r_rabbitpic[2477] <= 4'b1111;
        r_rabbitpic[2478] <= 4'b1111;
        r_rabbitpic[2479] <= 4'b1111;
        r_rabbitpic[2480] <= 4'b1111;
        r_rabbitpic[2481] <= 4'b1111;
        r_rabbitpic[2482] <= 4'b1111;
        r_rabbitpic[2483] <= 4'b1111;
        r_rabbitpic[2484] <= 4'b1111;
        r_rabbitpic[2485] <= 4'b1111;
        r_rabbitpic[2486] <= 4'b1111;
        r_rabbitpic[2487] <= 4'b1111;
        r_rabbitpic[2488] <= 4'b1111;
        r_rabbitpic[2489] <= 4'b1111;
        r_rabbitpic[2490] <= 4'b1111;
        r_rabbitpic[2491] <= 4'b1111;
        r_rabbitpic[2492] <= 4'b1111;
        r_rabbitpic[2493] <= 4'b1111;
        r_rabbitpic[2494] <= 4'b1111;
        r_rabbitpic[2495] <= 4'b1111;
        r_rabbitpic[2496] <= 4'b1111;
        r_rabbitpic[2497] <= 4'b1111;
        r_rabbitpic[2498] <= 4'b0000;
        r_rabbitpic[2499] <= 4'b0000;
        r_rabbitpic[2500] <= 4'b0000;
        r_rabbitpic[2501] <= 4'b0000;
        r_rabbitpic[2502] <= 4'b0000;
        r_rabbitpic[2503] <= 4'b0000;
        r_rabbitpic[2504] <= 4'b0000;
        r_rabbitpic[2505] <= 4'b0000;
        r_rabbitpic[2506] <= 4'b0000;
        r_rabbitpic[2507] <= 4'b0000;
        r_rabbitpic[2508] <= 4'b1111;
        r_rabbitpic[2509] <= 4'b1111;
        r_rabbitpic[2510] <= 4'b1111;
        r_rabbitpic[2511] <= 4'b0000;
        r_rabbitpic[2512] <= 4'b1111;
        r_rabbitpic[2513] <= 4'b1111;
        r_rabbitpic[2514] <= 4'b1111;
        r_rabbitpic[2515] <= 4'b0000;
        r_rabbitpic[2516] <= 4'b0000;
        r_rabbitpic[2517] <= 4'b1111;
        r_rabbitpic[2518] <= 4'b1111;
        r_rabbitpic[2519] <= 4'b0000;
        r_rabbitpic[2520] <= 4'b1111;
        r_rabbitpic[2521] <= 4'b1111;
        r_rabbitpic[2522] <= 4'b1111;
        r_rabbitpic[2523] <= 4'b1111;
        r_rabbitpic[2524] <= 4'b1111;
        r_rabbitpic[2525] <= 4'b1111;
        r_rabbitpic[2526] <= 4'b1111;
        r_rabbitpic[2527] <= 4'b1111;
        r_rabbitpic[2528] <= 4'b1111;
        r_rabbitpic[2529] <= 4'b1111;
        r_rabbitpic[2530] <= 4'b1111;
        r_rabbitpic[2531] <= 4'b1111;
        r_rabbitpic[2532] <= 4'b1111;
        r_rabbitpic[2533] <= 4'b1111;
        r_rabbitpic[2534] <= 4'b1111;
        r_rabbitpic[2535] <= 4'b1111;
        r_rabbitpic[2536] <= 4'b1111;
        r_rabbitpic[2537] <= 4'b1111;
        r_rabbitpic[2538] <= 4'b1111;
        r_rabbitpic[2539] <= 4'b1111;
        r_rabbitpic[2540] <= 4'b1111;
        r_rabbitpic[2541] <= 4'b1111;
        r_rabbitpic[2542] <= 4'b1111;
        r_rabbitpic[2543] <= 4'b1111;
        r_rabbitpic[2544] <= 4'b1111;
        r_rabbitpic[2545] <= 4'b1111;
        r_rabbitpic[2546] <= 4'b1111;
        r_rabbitpic[2547] <= 4'b1111;
        r_rabbitpic[2548] <= 4'b1111;
        r_rabbitpic[2549] <= 4'b0000;
        r_rabbitpic[2550] <= 4'b1111;
        r_rabbitpic[2551] <= 4'b1111;
        r_rabbitpic[2552] <= 4'b0000;
        r_rabbitpic[2553] <= 4'b0000;
        r_rabbitpic[2554] <= 4'b0000;
        r_rabbitpic[2555] <= 4'b1111;
        r_rabbitpic[2556] <= 4'b1111;
        r_rabbitpic[2557] <= 4'b1111;
        r_rabbitpic[2558] <= 4'b0000;
        r_rabbitpic[2559] <= 4'b0000;
        r_rabbitpic[2560] <= 4'b0000;
        r_rabbitpic[2561] <= 4'b0000;
        r_rabbitpic[2562] <= 4'b0000;
        r_rabbitpic[2563] <= 4'b0000;
        r_rabbitpic[2564] <= 4'b0000;
        r_rabbitpic[2565] <= 4'b0000;
        r_rabbitpic[2566] <= 4'b0000;
        r_rabbitpic[2567] <= 4'b1111;
        r_rabbitpic[2568] <= 4'b1111;
        r_rabbitpic[2569] <= 4'b1111;
        r_rabbitpic[2570] <= 4'b0000;
        r_rabbitpic[2571] <= 4'b0000;
        r_rabbitpic[2572] <= 4'b0000;
        r_rabbitpic[2573] <= 4'b0000;
        r_rabbitpic[2574] <= 4'b1111;
        r_rabbitpic[2575] <= 4'b1111;
        r_rabbitpic[2576] <= 4'b1111;
        r_rabbitpic[2577] <= 4'b1111;
        r_rabbitpic[2578] <= 4'b1111;
        r_rabbitpic[2579] <= 4'b1111;
        r_rabbitpic[2580] <= 4'b1111;
        r_rabbitpic[2581] <= 4'b1111;
        r_rabbitpic[2582] <= 4'b1111;
        r_rabbitpic[2583] <= 4'b1111;
        r_rabbitpic[2584] <= 4'b1111;
        r_rabbitpic[2585] <= 4'b1111;
        r_rabbitpic[2586] <= 4'b1111;
        r_rabbitpic[2587] <= 4'b1111;
        r_rabbitpic[2588] <= 4'b1111;
        r_rabbitpic[2589] <= 4'b1111;
        r_rabbitpic[2590] <= 4'b1111;
        r_rabbitpic[2591] <= 4'b1111;
        r_rabbitpic[2592] <= 4'b1111;
        r_rabbitpic[2593] <= 4'b1111;
        r_rabbitpic[2594] <= 4'b1111;
        r_rabbitpic[2595] <= 4'b1111;
        r_rabbitpic[2596] <= 4'b1111;
        r_rabbitpic[2597] <= 4'b1111;
        r_rabbitpic[2598] <= 4'b1111;
        r_rabbitpic[2599] <= 4'b1111;
        r_rabbitpic[2600] <= 4'b1111;
        r_rabbitpic[2601] <= 4'b1111;
        r_rabbitpic[2602] <= 4'b0000;
        r_rabbitpic[2603] <= 4'b0000;
        r_rabbitpic[2604] <= 4'b0000;
        r_rabbitpic[2605] <= 4'b1111;
        r_rabbitpic[2606] <= 4'b1111;
        r_rabbitpic[2607] <= 4'b0000;
        r_rabbitpic[2608] <= 4'b0000;
        r_rabbitpic[2609] <= 4'b1111;
        r_rabbitpic[2610] <= 4'b1111;
        r_rabbitpic[2611] <= 4'b1111;
        r_rabbitpic[2612] <= 4'b0000;
        r_rabbitpic[2613] <= 4'b0000;
        r_rabbitpic[2614] <= 4'b0000;
        r_rabbitpic[2615] <= 4'b1111;
        r_rabbitpic[2616] <= 4'b1111;
        r_rabbitpic[2617] <= 4'b1111;
        r_rabbitpic[2618] <= 4'b1111;
        r_rabbitpic[2619] <= 4'b1111;
        r_rabbitpic[2620] <= 4'b1111;
        r_rabbitpic[2621] <= 4'b1111;
        r_rabbitpic[2622] <= 4'b1111;
        r_rabbitpic[2623] <= 4'b1111;
        r_rabbitpic[2624] <= 4'b1111;
        r_rabbitpic[2625] <= 4'b0000;
        r_rabbitpic[2626] <= 4'b1111;
        r_rabbitpic[2627] <= 4'b1111;
        r_rabbitpic[2628] <= 4'b1111;
        r_rabbitpic[2629] <= 4'b1111;
        r_rabbitpic[2630] <= 4'b1111;
        r_rabbitpic[2631] <= 4'b1111;
        r_rabbitpic[2632] <= 4'b1111;
        r_rabbitpic[2633] <= 4'b1111;
        r_rabbitpic[2634] <= 4'b1111;
        r_rabbitpic[2635] <= 4'b1111;
        r_rabbitpic[2636] <= 4'b1111;
        r_rabbitpic[2637] <= 4'b1111;
        r_rabbitpic[2638] <= 4'b1111;
        r_rabbitpic[2639] <= 4'b1111;
        r_rabbitpic[2640] <= 4'b1111;
        r_rabbitpic[2641] <= 4'b1111;
        r_rabbitpic[2642] <= 4'b1111;
        r_rabbitpic[2643] <= 4'b1111;
        r_rabbitpic[2644] <= 4'b1111;
        r_rabbitpic[2645] <= 4'b1111;
        r_rabbitpic[2646] <= 4'b1111;
        r_rabbitpic[2647] <= 4'b1111;
        r_rabbitpic[2648] <= 4'b1111;
        r_rabbitpic[2649] <= 4'b1111;
        r_rabbitpic[2650] <= 4'b1111;
        r_rabbitpic[2651] <= 4'b1111;
        r_rabbitpic[2652] <= 4'b1111;
        r_rabbitpic[2653] <= 4'b1111;
        r_rabbitpic[2654] <= 4'b1111;
        r_rabbitpic[2655] <= 4'b1111;
        r_rabbitpic[2656] <= 4'b0000;
        r_rabbitpic[2657] <= 4'b1111;
        r_rabbitpic[2658] <= 4'b0000;
        r_rabbitpic[2659] <= 4'b1111;
        r_rabbitpic[2660] <= 4'b1111;
        r_rabbitpic[2661] <= 4'b0000;
        r_rabbitpic[2662] <= 4'b0000;
        r_rabbitpic[2663] <= 4'b1111;
        r_rabbitpic[2664] <= 4'b0000;
        r_rabbitpic[2665] <= 4'b1111;
        r_rabbitpic[2666] <= 4'b1111;
        r_rabbitpic[2667] <= 4'b0000;
        r_rabbitpic[2668] <= 4'b0000;
        r_rabbitpic[2669] <= 4'b0000;
        r_rabbitpic[2670] <= 4'b0000;
        r_rabbitpic[2671] <= 4'b0000;
        r_rabbitpic[2672] <= 4'b0000;
        r_rabbitpic[2673] <= 4'b0000;
        r_rabbitpic[2674] <= 4'b0000;
        r_rabbitpic[2675] <= 4'b0000;
        r_rabbitpic[2676] <= 4'b0000;
        r_rabbitpic[2677] <= 4'b0000;
        r_rabbitpic[2678] <= 4'b0000;
        r_rabbitpic[2679] <= 4'b0000;
        r_rabbitpic[2680] <= 4'b0000;
        r_rabbitpic[2681] <= 4'b1111;
        r_rabbitpic[2682] <= 4'b1111;
        r_rabbitpic[2683] <= 4'b1111;
        r_rabbitpic[2684] <= 4'b1111;
        r_rabbitpic[2685] <= 4'b1111;
        r_rabbitpic[2686] <= 4'b1111;
        r_rabbitpic[2687] <= 4'b1111;
        r_rabbitpic[2688] <= 4'b1111;
        r_rabbitpic[2689] <= 4'b1111;
        r_rabbitpic[2690] <= 4'b1111;
        r_rabbitpic[2691] <= 4'b1111;
        r_rabbitpic[2692] <= 4'b1111;
        r_rabbitpic[2693] <= 4'b1111;
        r_rabbitpic[2694] <= 4'b1111;
        r_rabbitpic[2695] <= 4'b1111;
        r_rabbitpic[2696] <= 4'b1111;
        r_rabbitpic[2697] <= 4'b1111;
        r_rabbitpic[2698] <= 4'b1111;
        r_rabbitpic[2699] <= 4'b1111;
        r_rabbitpic[2700] <= 4'b1111;
        r_rabbitpic[2701] <= 4'b1111;
        r_rabbitpic[2702] <= 4'b1111;
        r_rabbitpic[2703] <= 4'b1111;
        r_rabbitpic[2704] <= 4'b1111;
        r_rabbitpic[2705] <= 4'b1111;
        r_rabbitpic[2706] <= 4'b1111;
        r_rabbitpic[2707] <= 4'b1111;
        r_rabbitpic[2708] <= 4'b1111;
        r_rabbitpic[2709] <= 4'b1111;
        r_rabbitpic[2710] <= 4'b1111;
        r_rabbitpic[2711] <= 4'b0000;
        r_rabbitpic[2712] <= 4'b0000;
        r_rabbitpic[2713] <= 4'b1111;
        r_rabbitpic[2714] <= 4'b0000;
        r_rabbitpic[2715] <= 4'b0000;
        r_rabbitpic[2716] <= 4'b0000;
        r_rabbitpic[2717] <= 4'b1111;
        r_rabbitpic[2718] <= 4'b1111;
        r_rabbitpic[2719] <= 4'b1111;
        r_rabbitpic[2720] <= 4'b1111;
        r_rabbitpic[2721] <= 4'b1111;
        r_rabbitpic[2722] <= 4'b1111;
        r_rabbitpic[2723] <= 4'b1111;
        r_rabbitpic[2724] <= 4'b1111;
        r_rabbitpic[2725] <= 4'b1111;
        r_rabbitpic[2726] <= 4'b1111;
        r_rabbitpic[2727] <= 4'b1111;
        r_rabbitpic[2728] <= 4'b1111;
        r_rabbitpic[2729] <= 4'b1111;
        r_rabbitpic[2730] <= 4'b1111;
        r_rabbitpic[2731] <= 4'b1111;
        r_rabbitpic[2732] <= 4'b1111;
        r_rabbitpic[2733] <= 4'b1111;
        r_rabbitpic[2734] <= 4'b1111;
        r_rabbitpic[2735] <= 4'b1111;
        r_rabbitpic[2736] <= 4'b1111;
        r_rabbitpic[2737] <= 4'b1111;
        r_rabbitpic[2738] <= 4'b1111;
        r_rabbitpic[2739] <= 4'b1111;
        r_rabbitpic[2740] <= 4'b1111;
        r_rabbitpic[2741] <= 4'b1111;
        r_rabbitpic[2742] <= 4'b1111;
        r_rabbitpic[2743] <= 4'b1111;
        r_rabbitpic[2744] <= 4'b1111;
        r_rabbitpic[2745] <= 4'b1111;
        r_rabbitpic[2746] <= 4'b1111;
        r_rabbitpic[2747] <= 4'b1111;
        r_rabbitpic[2748] <= 4'b1111;
        r_rabbitpic[2749] <= 4'b1111;
        r_rabbitpic[2750] <= 4'b1111;
        r_rabbitpic[2751] <= 4'b1111;
        r_rabbitpic[2752] <= 4'b1111;
        r_rabbitpic[2753] <= 4'b1111;
        r_rabbitpic[2754] <= 4'b1111;
        r_rabbitpic[2755] <= 4'b1111;
        r_rabbitpic[2756] <= 4'b1111;
        r_rabbitpic[2757] <= 4'b1111;
        r_rabbitpic[2758] <= 4'b1111;
        r_rabbitpic[2759] <= 4'b1111;
        r_rabbitpic[2760] <= 4'b1111;
        r_rabbitpic[2761] <= 4'b1111;
        r_rabbitpic[2762] <= 4'b1111;
        r_rabbitpic[2763] <= 4'b1111;
        r_rabbitpic[2764] <= 4'b1111;
        r_rabbitpic[2765] <= 4'b1111;
        r_rabbitpic[2766] <= 4'b1111;
        r_rabbitpic[2767] <= 4'b0000;
        r_rabbitpic[2768] <= 4'b0000;
        r_rabbitpic[2769] <= 4'b1111;
        r_rabbitpic[2770] <= 4'b1111;
        r_rabbitpic[2771] <= 4'b1111;
        r_rabbitpic[2772] <= 4'b1111;
        r_rabbitpic[2773] <= 4'b1111;
        r_rabbitpic[2774] <= 4'b1111;
        r_rabbitpic[2775] <= 4'b1111;
        r_rabbitpic[2776] <= 4'b1111;
        r_rabbitpic[2777] <= 4'b1111;
        r_rabbitpic[2778] <= 4'b1111;
        r_rabbitpic[2779] <= 4'b1111;
        r_rabbitpic[2780] <= 4'b1111;
        r_rabbitpic[2781] <= 4'b1111;
        r_rabbitpic[2782] <= 4'b1111;
        r_rabbitpic[2783] <= 4'b1111;
        r_rabbitpic[2784] <= 4'b1111;
        r_rabbitpic[2785] <= 4'b1111;
        r_rabbitpic[2786] <= 4'b1111;
        r_rabbitpic[2787] <= 4'b1111;
        r_rabbitpic[2788] <= 4'b1111;
        r_rabbitpic[2789] <= 4'b1111;
        r_rabbitpic[2790] <= 4'b1111;
        r_rabbitpic[2791] <= 4'b1111;
        r_rabbitpic[2792] <= 4'b1111;
        r_rabbitpic[2793] <= 4'b1111;
        r_rabbitpic[2794] <= 4'b1111;
        r_rabbitpic[2795] <= 4'b1111;
        r_rabbitpic[2796] <= 4'b1111;
        r_rabbitpic[2797] <= 4'b1111;
        r_rabbitpic[2798] <= 4'b1111;
        r_rabbitpic[2799] <= 4'b1111;
        r_rabbitpic[2800] <= 4'b1111;
        r_rabbitpic[2801] <= 4'b1111;
        r_rabbitpic[2802] <= 4'b1111;
        r_rabbitpic[2803] <= 4'b1111;
        r_rabbitpic[2804] <= 4'b1111;
        r_rabbitpic[2805] <= 4'b1111;
        r_rabbitpic[2806] <= 4'b1111;
        r_rabbitpic[2807] <= 4'b1111;
        r_rabbitpic[2808] <= 4'b1111;
        r_rabbitpic[2809] <= 4'b1111;
        r_rabbitpic[2810] <= 4'b1111;
        r_rabbitpic[2811] <= 4'b1111;
        r_rabbitpic[2812] <= 4'b1111;
        r_rabbitpic[2813] <= 4'b1111;
        r_rabbitpic[2814] <= 4'b1111;
        r_rabbitpic[2815] <= 4'b1111;
        r_rabbitpic[2816] <= 4'b1111;
        r_rabbitpic[2817] <= 4'b1111;
        r_rabbitpic[2818] <= 4'b1111;
        r_rabbitpic[2819] <= 4'b1111;
        r_rabbitpic[2820] <= 4'b1111;
        r_rabbitpic[2821] <= 4'b1111;
        r_rabbitpic[2822] <= 4'b1111;
        r_rabbitpic[2823] <= 4'b1111;
        r_rabbitpic[2824] <= 4'b1111;
        r_rabbitpic[2825] <= 4'b1111;
        r_rabbitpic[2826] <= 4'b1111;
        r_rabbitpic[2827] <= 4'b1111;
        r_rabbitpic[2828] <= 4'b1111;
        r_rabbitpic[2829] <= 4'b1111;
        r_rabbitpic[2830] <= 4'b1111;
        r_rabbitpic[2831] <= 4'b1111;
        r_rabbitpic[2832] <= 4'b1111;
        r_rabbitpic[2833] <= 4'b1111;
        r_rabbitpic[2834] <= 4'b1111;
        r_rabbitpic[2835] <= 4'b1111;
        r_rabbitpic[2836] <= 4'b1111;
        r_rabbitpic[2837] <= 4'b1111;
        r_rabbitpic[2838] <= 4'b1111;
        r_rabbitpic[2839] <= 4'b1111;
        r_rabbitpic[2840] <= 4'b1111;
        r_rabbitpic[2841] <= 4'b1111;
        r_rabbitpic[2842] <= 4'b1111;
        r_rabbitpic[2843] <= 4'b1111;
        r_rabbitpic[2844] <= 4'b1111;
        r_rabbitpic[2845] <= 4'b1111;
        r_rabbitpic[2846] <= 4'b1111;
        r_rabbitpic[2847] <= 4'b1111;
        r_rabbitpic[2848] <= 4'b1111;
        r_rabbitpic[2849] <= 4'b1111;
        r_rabbitpic[2850] <= 4'b1111;
        r_rabbitpic[2851] <= 4'b1111;
        r_rabbitpic[2852] <= 4'b1111;
        r_rabbitpic[2853] <= 4'b1111;
        r_rabbitpic[2854] <= 4'b1111;
        r_rabbitpic[2855] <= 4'b1111;
        r_rabbitpic[2856] <= 4'b1111;
        r_rabbitpic[2857] <= 4'b1111;
        r_rabbitpic[2858] <= 4'b1111;
        r_rabbitpic[2859] <= 4'b1111;
        r_rabbitpic[2860] <= 4'b1111;
        r_rabbitpic[2861] <= 4'b1111;
        r_rabbitpic[2862] <= 4'b1111;
        r_rabbitpic[2863] <= 4'b1111;
        r_rabbitpic[2864] <= 4'b1111;
        r_rabbitpic[2865] <= 4'b1111;
        r_rabbitpic[2866] <= 4'b1111;
        r_rabbitpic[2867] <= 4'b1111;
        r_rabbitpic[2868] <= 4'b1111;
        r_rabbitpic[2869] <= 4'b1111;
        r_rabbitpic[2870] <= 4'b1111;
        r_rabbitpic[2871] <= 4'b1111;
        r_rabbitpic[2872] <= 4'b1111;
        r_rabbitpic[2873] <= 4'b1111;
        r_rabbitpic[2874] <= 4'b1111;
        r_rabbitpic[2875] <= 4'b1111;
        r_rabbitpic[2876] <= 4'b1111;
        r_rabbitpic[2877] <= 4'b1111;
        r_rabbitpic[2878] <= 4'b1111;
        r_rabbitpic[2879] <= 4'b1111;
        r_rabbitpic[2880] <= 4'b1111;
        r_rabbitpic[2881] <= 4'b1111;
        r_rabbitpic[2882] <= 4'b1111;
        r_rabbitpic[2883] <= 4'b1111;
        r_rabbitpic[2884] <= 4'b1111;
        r_rabbitpic[2885] <= 4'b1111;
        r_rabbitpic[2886] <= 4'b1111;
        r_rabbitpic[2887] <= 4'b1111;
        r_rabbitpic[2888] <= 4'b1111;
        r_rabbitpic[2889] <= 4'b1111;
        r_rabbitpic[2890] <= 4'b1111;
        r_rabbitpic[2891] <= 4'b1111;
        r_rabbitpic[2892] <= 4'b1111;
        r_rabbitpic[2893] <= 4'b1111;
        r_rabbitpic[2894] <= 4'b1111;
        r_rabbitpic[2895] <= 4'b1111;
        r_rabbitpic[2896] <= 4'b1111;
        r_rabbitpic[2897] <= 4'b1111;
        r_rabbitpic[2898] <= 4'b1111;
        r_rabbitpic[2899] <= 4'b1111;
        r_rabbitpic[2900] <= 4'b1111;
        r_rabbitpic[2901] <= 4'b1111;
        r_rabbitpic[2902] <= 4'b1111;
        r_rabbitpic[2903] <= 4'b1111;
        r_rabbitpic[2904] <= 4'b1111;
        r_rabbitpic[2905] <= 4'b1111;
        r_rabbitpic[2906] <= 4'b1111;
        r_rabbitpic[2907] <= 4'b1111;
        r_rabbitpic[2908] <= 4'b1111;
        r_rabbitpic[2909] <= 4'b1111;
        r_rabbitpic[2910] <= 4'b1111;
        r_rabbitpic[2911] <= 4'b1111;
        r_rabbitpic[2912] <= 4'b1111;
        r_rabbitpic[2913] <= 4'b1111;
        r_rabbitpic[2914] <= 4'b1111;
        r_rabbitpic[2915] <= 4'b1111;
        r_rabbitpic[2916] <= 4'b1111;
        r_rabbitpic[2917] <= 4'b1111;
        r_rabbitpic[2918] <= 4'b1111;
        r_rabbitpic[2919] <= 4'b1111;
        r_rabbitpic[2920] <= 4'b1111;
        r_rabbitpic[2921] <= 4'b1111;
        r_rabbitpic[2922] <= 4'b1111;
        r_rabbitpic[2923] <= 4'b1111;
        r_rabbitpic[2924] <= 4'b1111;
        r_rabbitpic[2925] <= 4'b1111;
        r_rabbitpic[2926] <= 4'b1111;
        r_rabbitpic[2927] <= 4'b1111;
        r_rabbitpic[2928] <= 4'b1111;
        r_rabbitpic[2929] <= 4'b1111;
        r_rabbitpic[2930] <= 4'b1111;
        r_rabbitpic[2931] <= 4'b1111;
        r_rabbitpic[2932] <= 4'b1111;
        r_rabbitpic[2933] <= 4'b1111;
        r_rabbitpic[2934] <= 4'b1111;
        r_rabbitpic[2935] <= 4'b1111;
        r_rabbitpic[2936] <= 4'b1111;
        r_rabbitpic[2937] <= 4'b1111;
        r_rabbitpic[2938] <= 4'b1111;
        r_rabbitpic[2939] <= 4'b1111;
        r_rabbitpic[2940] <= 4'b1111;
        r_rabbitpic[2941] <= 4'b1111;
        r_rabbitpic[2942] <= 4'b1111;
        r_rabbitpic[2943] <= 4'b1111;
        r_rabbitpic[2944] <= 4'b1111;
        r_rabbitpic[2945] <= 4'b1111;
        r_rabbitpic[2946] <= 4'b1111;
        r_rabbitpic[2947] <= 4'b1111;
        r_rabbitpic[2948] <= 4'b1111;
        r_rabbitpic[2949] <= 4'b1111;
        r_rabbitpic[2950] <= 4'b1111;
        r_rabbitpic[2951] <= 4'b1111;
        r_rabbitpic[2952] <= 4'b1111;
        r_rabbitpic[2953] <= 4'b1111;
        r_rabbitpic[2954] <= 4'b1111;
        r_rabbitpic[2955] <= 4'b1111;
        r_rabbitpic[2956] <= 4'b1111;
        r_rabbitpic[2957] <= 4'b1111;
        r_rabbitpic[2958] <= 4'b1111;
        r_rabbitpic[2959] <= 4'b1111;
        r_rabbitpic[2960] <= 4'b1111;
        r_rabbitpic[2961] <= 4'b1111;
        r_rabbitpic[2962] <= 4'b1111;
        r_rabbitpic[2963] <= 4'b1111;
        r_rabbitpic[2964] <= 4'b1111;
        r_rabbitpic[2965] <= 4'b1111;
        r_rabbitpic[2966] <= 4'b1111;
        r_rabbitpic[2967] <= 4'b1111;
        r_rabbitpic[2968] <= 4'b1111;
        r_rabbitpic[2969] <= 4'b1111;
        r_rabbitpic[2970] <= 4'b1111;
        r_rabbitpic[2971] <= 4'b1111;
        r_rabbitpic[2972] <= 4'b1111;
        r_rabbitpic[2973] <= 4'b1111;
        r_rabbitpic[2974] <= 4'b1111;
        r_rabbitpic[2975] <= 4'b1111;
        r_rabbitpic[2976] <= 4'b1111;
        r_rabbitpic[2977] <= 4'b1111;
        r_rabbitpic[2978] <= 4'b1111;
        r_rabbitpic[2979] <= 4'b1111;
        r_rabbitpic[2980] <= 4'b1111;
        r_rabbitpic[2981] <= 4'b1111;
        r_rabbitpic[2982] <= 4'b1111;
        r_rabbitpic[2983] <= 4'b1111;
        r_rabbitpic[2984] <= 4'b1111;
        r_rabbitpic[2985] <= 4'b1111;
        r_rabbitpic[2986] <= 4'b1111;
        r_rabbitpic[2987] <= 4'b1111;
        r_rabbitpic[2988] <= 4'b1111;
        r_rabbitpic[2989] <= 4'b1111;
        r_rabbitpic[2990] <= 4'b1111;
        r_rabbitpic[2991] <= 4'b1111;
        r_rabbitpic[2992] <= 4'b1111;
        r_rabbitpic[2993] <= 4'b1111;
        r_rabbitpic[2994] <= 4'b1111;
        r_rabbitpic[2995] <= 4'b1111;
        r_rabbitpic[2996] <= 4'b1111;
        r_rabbitpic[2997] <= 4'b1111;
        r_rabbitpic[2998] <= 4'b1111;
        r_rabbitpic[2999] <= 4'b1111;
        r_rabbitpic[3000] <= 4'b1111;
        r_rabbitpic[3001] <= 4'b1111;
        r_rabbitpic[3002] <= 4'b1111;
        r_rabbitpic[3003] <= 4'b1111;
        r_rabbitpic[3004] <= 4'b1111;
        r_rabbitpic[3005] <= 4'b1111;
        r_rabbitpic[3006] <= 4'b1111;
        r_rabbitpic[3007] <= 4'b1111;
        r_rabbitpic[3008] <= 4'b1111;
        r_rabbitpic[3009] <= 4'b1111;
        r_rabbitpic[3010] <= 4'b1111;
        r_rabbitpic[3011] <= 4'b1111;
        r_rabbitpic[3012] <= 4'b1111;
        r_rabbitpic[3013] <= 4'b1111;
        r_rabbitpic[3014] <= 4'b1111;
        r_rabbitpic[3015] <= 4'b1111;
        r_rabbitpic[3016] <= 4'b1111;
        r_rabbitpic[3017] <= 4'b1111;
        r_rabbitpic[3018] <= 4'b1111;
        r_rabbitpic[3019] <= 4'b1111;
        r_rabbitpic[3020] <= 4'b1111;
        r_rabbitpic[3021] <= 4'b1111;
        r_rabbitpic[3022] <= 4'b1111;
        r_rabbitpic[3023] <= 4'b1111;
        r_rabbitpic[3024] <= 4'b1111;

    end
endmodule

   